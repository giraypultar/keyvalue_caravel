magic
tech sky130A
magscale 1 2
timestamp 1641005295
<< locali >>
rect 568957 525351 568991 540345
rect 568957 495363 568991 503013
rect 568957 485095 568991 486421
rect 567761 69411 567795 69785
rect 567669 69207 567703 69377
rect 69029 68731 69063 68969
rect 72617 68323 72651 68493
rect 79333 67643 79367 67949
rect 152105 67643 152139 68629
rect 154313 67643 154347 68765
rect 178049 67847 178083 68901
rect 182189 67847 182223 68833
rect 186053 67847 186087 68833
rect 190377 67847 190411 68901
rect 197369 68255 197403 68969
rect 200037 68255 200071 68969
rect 81541 64991 81575 66045
rect 73997 3451 74031 3553
rect 94973 3383 95007 3553
<< viali >>
rect 568957 540345 568991 540379
rect 568957 525317 568991 525351
rect 568957 503013 568991 503047
rect 568957 495329 568991 495363
rect 568957 486421 568991 486455
rect 568957 485061 568991 485095
rect 567761 69785 567795 69819
rect 567669 69377 567703 69411
rect 567761 69377 567795 69411
rect 567669 69173 567703 69207
rect 69029 68969 69063 69003
rect 197369 68969 197403 69003
rect 178049 68901 178083 68935
rect 69029 68697 69063 68731
rect 154313 68765 154347 68799
rect 152105 68629 152139 68663
rect 72617 68493 72651 68527
rect 72617 68289 72651 68323
rect 79333 67949 79367 67983
rect 79333 67609 79367 67643
rect 152105 67609 152139 67643
rect 190377 68901 190411 68935
rect 178049 67813 178083 67847
rect 182189 68833 182223 68867
rect 182189 67813 182223 67847
rect 186053 68833 186087 68867
rect 186053 67813 186087 67847
rect 197369 68221 197403 68255
rect 200037 68969 200071 69003
rect 200037 68221 200071 68255
rect 190377 67813 190411 67847
rect 154313 67609 154347 67643
rect 81541 66045 81575 66079
rect 81541 64957 81575 64991
rect 73997 3553 74031 3587
rect 73997 3417 74031 3451
rect 94973 3553 95007 3587
rect 94973 3349 95007 3383
<< metal1 >>
rect 283834 700816 283840 700868
rect 283892 700856 283898 700868
rect 439590 700856 439596 700868
rect 283892 700828 439596 700856
rect 283892 700816 283898 700828
rect 439590 700816 439596 700828
rect 439648 700816 439654 700868
rect 318702 700748 318708 700800
rect 318760 700788 318766 700800
rect 478506 700788 478512 700800
rect 318760 700760 478512 700788
rect 318760 700748 318766 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 170306 700680 170312 700732
rect 170364 700720 170370 700732
rect 333974 700720 333980 700732
rect 170364 700692 333980 700720
rect 170364 700680 170370 700692
rect 333974 700680 333980 700692
rect 334032 700680 334038 700732
rect 348786 700680 348792 700732
rect 348844 700720 348850 700732
rect 439498 700720 439504 700732
rect 348844 700692 439504 700720
rect 348844 700680 348850 700692
rect 439498 700680 439504 700692
rect 439556 700680 439562 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 418154 700652 418160 700664
rect 154172 700624 418160 700652
rect 154172 700612 154178 700624
rect 418154 700612 418160 700624
rect 418212 700612 418218 700664
rect 300118 700544 300124 700596
rect 300176 700584 300182 700596
rect 570322 700584 570328 700596
rect 300176 700556 570328 700584
rect 300176 700544 300182 700556
rect 570322 700544 570328 700556
rect 570380 700544 570386 700596
rect 277302 700476 277308 700528
rect 277360 700516 277366 700528
rect 559650 700516 559656 700528
rect 277360 700488 559656 700516
rect 277360 700476 277366 700488
rect 559650 700476 559656 700488
rect 559708 700476 559714 700528
rect 69842 700408 69848 700460
rect 69900 700448 69906 700460
rect 364978 700448 364984 700460
rect 69900 700420 364984 700448
rect 69900 700408 69906 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 413646 700408 413652 700460
rect 413704 700448 413710 700460
rect 568850 700448 568856 700460
rect 413704 700420 568856 700448
rect 413704 700408 413710 700420
rect 568850 700408 568856 700420
rect 568908 700408 568914 700460
rect 89162 700340 89168 700392
rect 89220 700380 89226 700392
rect 424318 700380 424324 700392
rect 89220 700352 424324 700380
rect 89220 700340 89226 700352
rect 424318 700340 424324 700352
rect 424376 700340 424382 700392
rect 543458 700340 543464 700392
rect 543516 700380 543522 700392
rect 568574 700380 568580 700392
rect 543516 700352 568580 700380
rect 543516 700340 543522 700352
rect 568574 700340 568580 700352
rect 568632 700340 568638 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 105538 700312 105544 700324
rect 40552 700284 105544 700312
rect 40552 700272 40558 700284
rect 105538 700272 105544 700284
rect 105596 700272 105602 700324
rect 218974 700272 218980 700324
rect 219032 700312 219038 700324
rect 570046 700312 570052 700324
rect 219032 700284 570052 700312
rect 219032 700272 219038 700284
rect 570046 700272 570052 700284
rect 570104 700272 570110 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 494790 699660 494796 699712
rect 494848 699700 494854 699712
rect 495342 699700 495348 699712
rect 494848 699672 495348 699700
rect 494848 699660 494854 699672
rect 495342 699660 495348 699672
rect 495400 699660 495406 699712
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 569954 683176 569960 683188
rect 3476 683148 569960 683176
rect 3476 683136 3482 683148
rect 569954 683136 569960 683148
rect 570012 683136 570018 683188
rect 576210 683136 576216 683188
rect 576268 683176 576274 683188
rect 580166 683176 580172 683188
rect 576268 683148 580172 683176
rect 576268 683136 576274 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 2774 671032 2780 671084
rect 2832 671072 2838 671084
rect 4798 671072 4804 671084
rect 2832 671044 4804 671072
rect 2832 671032 2838 671044
rect 4798 671032 4804 671044
rect 4856 671032 4862 671084
rect 573358 670692 573364 670744
rect 573416 670732 573422 670744
rect 580166 670732 580172 670744
rect 573416 670704 580172 670732
rect 573416 670692 573422 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 570414 632108 570420 632120
rect 3476 632080 570420 632108
rect 3476 632068 3482 632080
rect 570414 632068 570420 632080
rect 570472 632068 570478 632120
rect 68738 630640 68744 630692
rect 68796 630680 68802 630692
rect 580166 630680 580172 630692
rect 68796 630652 580172 630680
rect 68796 630640 68802 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 256602 616836 256608 616888
rect 256660 616876 256666 616888
rect 580166 616876 580172 616888
rect 256660 616848 580172 616876
rect 256660 616836 256666 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 2774 579912 2780 579964
rect 2832 579952 2838 579964
rect 4890 579952 4896 579964
rect 2832 579924 4896 579952
rect 2832 579912 2838 579924
rect 4890 579912 4896 579924
rect 4948 579912 4954 579964
rect 574738 576852 574744 576904
rect 574796 576892 574802 576904
rect 580166 576892 580172 576904
rect 574796 576864 580172 576892
rect 574796 576852 574802 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 105538 571276 105544 571328
rect 105596 571316 105602 571328
rect 107194 571316 107200 571328
rect 105596 571288 107200 571316
rect 105596 571276 105602 571288
rect 107194 571276 107200 571288
rect 107252 571276 107258 571328
rect 276474 571276 276480 571328
rect 276532 571316 276538 571328
rect 277302 571316 277308 571328
rect 276532 571288 277308 571316
rect 276532 571276 276538 571288
rect 277302 571276 277308 571288
rect 277360 571276 277366 571328
rect 64138 571004 64144 571056
rect 64196 571044 64202 571056
rect 186498 571044 186504 571056
rect 64196 571016 186504 571044
rect 64196 571004 64202 571016
rect 186498 571004 186504 571016
rect 186556 571004 186562 571056
rect 10318 570936 10324 570988
rect 10376 570976 10382 570988
rect 530210 570976 530216 570988
rect 10376 570948 530216 570976
rect 10376 570936 10382 570948
rect 530210 570936 530216 570948
rect 530268 570936 530274 570988
rect 58618 570800 58624 570852
rect 58676 570840 58682 570852
rect 138842 570840 138848 570852
rect 58676 570812 138848 570840
rect 58676 570800 58682 570812
rect 138842 570800 138848 570812
rect 138900 570800 138906 570852
rect 57238 570732 57244 570784
rect 57296 570772 57302 570784
rect 149514 570772 149520 570784
rect 57296 570744 149520 570772
rect 57296 570732 57302 570744
rect 149514 570732 149520 570744
rect 149572 570732 149578 570784
rect 255314 570732 255320 570784
rect 255372 570772 255378 570784
rect 256602 570772 256608 570784
rect 255372 570744 256608 570772
rect 255372 570732 255378 570744
rect 256602 570732 256608 570744
rect 256660 570732 256666 570784
rect 439498 570732 439504 570784
rect 439556 570772 439562 570784
rect 472066 570772 472072 570784
rect 439556 570744 472072 570772
rect 439556 570732 439562 570744
rect 472066 570732 472072 570744
rect 472124 570732 472130 570784
rect 495342 570732 495348 570784
rect 495400 570772 495406 570784
rect 535546 570772 535552 570784
rect 495400 570744 535552 570772
rect 495400 570732 495406 570744
rect 535546 570732 535552 570744
rect 535604 570732 535610 570784
rect 54478 570664 54484 570716
rect 54536 570704 54542 570716
rect 165338 570704 165344 570716
rect 54536 570676 165344 570704
rect 54536 570664 54542 570676
rect 165338 570664 165344 570676
rect 165396 570664 165402 570716
rect 439590 570664 439596 570716
rect 439648 570704 439654 570716
rect 556706 570704 556712 570716
rect 439648 570676 556712 570704
rect 439648 570664 439654 570676
rect 556706 570664 556712 570676
rect 556764 570664 556770 570716
rect 12342 570596 12348 570648
rect 12400 570636 12406 570648
rect 123018 570636 123024 570648
rect 12400 570608 123024 570636
rect 12400 570596 12406 570608
rect 123018 570596 123024 570608
rect 123076 570596 123082 570648
rect 424318 570596 424324 570648
rect 424376 570636 424382 570648
rect 561858 570636 561864 570648
rect 424376 570608 561864 570636
rect 424376 570596 424382 570608
rect 561858 570596 561864 570608
rect 561916 570596 561922 570648
rect 65518 570528 65524 570580
rect 65576 570568 65582 570580
rect 191834 570568 191840 570580
rect 65576 570540 191840 570568
rect 65576 570528 65582 570540
rect 191834 570528 191840 570540
rect 191892 570528 191898 570580
rect 68830 570460 68836 570512
rect 68888 570500 68894 570512
rect 239306 570500 239312 570512
rect 68888 570472 239312 570500
rect 68888 570460 68894 570472
rect 239306 570460 239312 570472
rect 239364 570460 239370 570512
rect 22738 570392 22744 570444
rect 22796 570432 22802 570444
rect 196986 570432 196992 570444
rect 22796 570404 196992 570432
rect 22796 570392 22802 570404
rect 196986 570392 196992 570404
rect 197044 570392 197050 570444
rect 178126 570324 178132 570376
rect 178184 570364 178190 570376
rect 456242 570364 456248 570376
rect 178184 570336 456248 570364
rect 178184 570324 178190 570336
rect 456242 570324 456248 570336
rect 456300 570324 456306 570376
rect 39298 570256 39304 570308
rect 39356 570296 39362 570308
rect 350442 570296 350448 570308
rect 39356 570268 350448 570296
rect 39356 570256 39362 570268
rect 350442 570256 350448 570268
rect 350500 570256 350506 570308
rect 408586 570256 408592 570308
rect 408644 570296 408650 570308
rect 569310 570296 569316 570308
rect 408644 570268 569316 570296
rect 408644 570256 408650 570268
rect 569310 570256 569316 570268
rect 569368 570256 569374 570308
rect 50338 570188 50344 570240
rect 50396 570228 50402 570240
rect 450906 570228 450912 570240
rect 50396 570200 450912 570228
rect 50396 570188 50402 570200
rect 450906 570188 450912 570200
rect 450964 570188 450970 570240
rect 69658 570120 69664 570172
rect 69716 570160 69722 570172
rect 477402 570160 477408 570172
rect 69716 570132 477408 570160
rect 69716 570120 69722 570132
rect 477402 570120 477408 570132
rect 477460 570120 477466 570172
rect 66070 570052 66076 570104
rect 66128 570092 66134 570104
rect 487890 570092 487896 570104
rect 66128 570064 487896 570092
rect 66128 570052 66134 570064
rect 487890 570052 487896 570064
rect 487948 570052 487954 570104
rect 26878 569984 26884 570036
rect 26936 570024 26942 570036
rect 509050 570024 509056 570036
rect 26936 569996 509056 570024
rect 26936 569984 26942 569996
rect 509050 569984 509056 569996
rect 509108 569984 509114 570036
rect 68922 569916 68928 569968
rect 68980 569956 68986 569968
rect 75362 569956 75368 569968
rect 68980 569928 75368 569956
rect 68980 569916 68986 569928
rect 75362 569916 75368 569928
rect 75420 569916 75426 569968
rect 234154 568216 234160 568268
rect 234212 568256 234218 568268
rect 573450 568256 573456 568268
rect 234212 568228 573456 568256
rect 234212 568216 234218 568228
rect 573450 568216 573456 568228
rect 573508 568216 573514 568268
rect 11698 568148 11704 568200
rect 11756 568188 11762 568200
rect 355778 568188 355784 568200
rect 11756 568160 355784 568188
rect 11756 568148 11762 568160
rect 355778 568148 355784 568160
rect 355836 568148 355842 568200
rect 10410 568080 10416 568132
rect 10468 568120 10474 568132
rect 360930 568120 360936 568132
rect 10468 568092 360936 568120
rect 10468 568080 10474 568092
rect 360930 568080 360936 568092
rect 360988 568080 360994 568132
rect 398098 568080 398104 568132
rect 398156 568120 398162 568132
rect 576302 568120 576308 568132
rect 398156 568092 576308 568120
rect 398156 568080 398162 568092
rect 576302 568080 576308 568092
rect 576360 568080 576366 568132
rect 5074 568012 5080 568064
rect 5132 568052 5138 568064
rect 218330 568052 218336 568064
rect 5132 568024 218336 568052
rect 5132 568012 5138 568024
rect 218330 568012 218336 568024
rect 218388 568012 218394 568064
rect 223298 568012 223304 568064
rect 223356 568052 223362 568064
rect 580258 568052 580264 568064
rect 223356 568024 580264 568052
rect 223356 568012 223362 568024
rect 580258 568012 580264 568024
rect 580316 568012 580322 568064
rect 7650 567944 7656 567996
rect 7708 567984 7714 567996
rect 365990 567984 365996 567996
rect 7708 567956 365996 567984
rect 7708 567944 7714 567956
rect 365990 567944 365996 567956
rect 366048 567944 366054 567996
rect 371970 567944 371976 567996
rect 372028 567984 372034 567996
rect 577498 567984 577504 567996
rect 372028 567956 577504 567984
rect 372028 567944 372034 567956
rect 577498 567944 577504 567956
rect 577556 567944 577562 567996
rect 208026 567876 208032 567928
rect 208084 567916 208090 567928
rect 573542 567916 573548 567928
rect 208084 567888 573548 567916
rect 208084 567876 208090 567888
rect 573542 567876 573548 567888
rect 573600 567876 573606 567928
rect 46842 567808 46848 567860
rect 46900 567848 46906 567860
rect 424134 567848 424140 567860
rect 46900 567820 424140 567848
rect 46900 567808 46906 567820
rect 424134 567808 424140 567820
rect 424192 567808 424198 567860
rect 3418 567740 3424 567792
rect 3476 567780 3482 567792
rect 159726 567780 159732 567792
rect 3476 567752 159732 567780
rect 3476 567740 3482 567752
rect 159726 567740 159732 567752
rect 159784 567740 159790 567792
rect 202690 567740 202696 567792
rect 202748 567780 202754 567792
rect 580350 567780 580356 567792
rect 202748 567752 580356 567780
rect 202748 567740 202754 567752
rect 580350 567740 580356 567752
rect 580408 567740 580414 567792
rect 44082 567672 44088 567724
rect 44140 567712 44146 567724
rect 429470 567712 429476 567724
rect 44140 567684 429476 567712
rect 44140 567672 44146 567684
rect 429470 567672 429476 567684
rect 429528 567672 429534 567724
rect 11790 567604 11796 567656
rect 11848 567644 11854 567656
rect 434806 567644 434812 567656
rect 11848 567616 434812 567644
rect 11848 567604 11854 567616
rect 434806 567604 434812 567616
rect 434864 567604 434870 567656
rect 445754 567604 445760 567656
rect 445812 567644 445818 567656
rect 574922 567644 574928 567656
rect 445812 567616 574928 567644
rect 445812 567604 445818 567616
rect 574922 567604 574928 567616
rect 574980 567604 574986 567656
rect 62022 567536 62028 567588
rect 62080 567576 62086 567588
rect 492950 567576 492956 567588
rect 62080 567548 492956 567576
rect 62080 567536 62086 567548
rect 492950 567536 492956 567548
rect 493008 567536 493014 567588
rect 118050 567468 118056 567520
rect 118108 567508 118114 567520
rect 574830 567508 574836 567520
rect 118108 567480 574836 567508
rect 118108 567468 118114 567480
rect 574830 567468 574836 567480
rect 574888 567468 574894 567520
rect 112806 567400 112812 567452
rect 112864 567440 112870 567452
rect 576118 567440 576124 567452
rect 112864 567412 576124 567440
rect 112864 567400 112870 567412
rect 576118 567400 576124 567412
rect 576176 567400 576182 567452
rect 39390 567332 39396 567384
rect 39448 567372 39454 567384
rect 514110 567372 514116 567384
rect 39448 567344 514116 567372
rect 39448 567332 39454 567344
rect 514110 567332 514116 567344
rect 514168 567332 514174 567384
rect 66162 567264 66168 567316
rect 66220 567304 66226 567316
rect 69934 567304 69940 567316
rect 66220 567276 69940 567304
rect 66220 567264 66226 567276
rect 69934 567264 69940 567276
rect 69992 567264 69998 567316
rect 91738 567264 91744 567316
rect 91796 567304 91802 567316
rect 91796 567276 93854 567304
rect 91796 567264 91802 567276
rect 93826 567236 93854 567276
rect 96706 567264 96712 567316
rect 96764 567304 96770 567316
rect 571242 567304 571248 567316
rect 96764 567276 571248 567304
rect 96764 567264 96770 567276
rect 571242 567264 571248 567276
rect 571300 567264 571306 567316
rect 570598 567236 570604 567248
rect 93826 567208 570604 567236
rect 570598 567196 570604 567208
rect 570656 567196 570662 567248
rect 3602 566448 3608 566500
rect 3660 566488 3666 566500
rect 570230 566488 570236 566500
rect 3660 566460 570236 566488
rect 3660 566448 3666 566460
rect 570230 566448 570236 566460
rect 570288 566448 570294 566500
rect 3510 566312 3516 566364
rect 3568 566352 3574 566364
rect 7558 566352 7564 566364
rect 3568 566324 7564 566352
rect 3568 566312 3574 566324
rect 7558 566312 7564 566324
rect 7616 566312 7622 566364
rect 568758 566012 568764 566024
rect 567166 565984 568764 566012
rect 567166 565944 567194 565984
rect 568758 565972 568764 565984
rect 568816 565972 568822 566024
rect 547846 565916 567194 565944
rect 69014 565836 69020 565888
rect 69072 565876 69078 565888
rect 547846 565876 547874 565916
rect 568574 565904 568580 565956
rect 568632 565944 568638 565956
rect 569402 565944 569408 565956
rect 568632 565916 569408 565944
rect 568632 565904 568638 565916
rect 569402 565904 569408 565916
rect 569460 565904 569466 565956
rect 69072 565848 547874 565876
rect 69072 565836 69078 565848
rect 571242 564340 571248 564392
rect 571300 564380 571306 564392
rect 580166 564380 580172 564392
rect 571300 564352 580172 564380
rect 571300 564340 571306 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 68646 561688 68652 561740
rect 68704 561728 68710 561740
rect 69014 561728 69020 561740
rect 68704 561700 69020 561728
rect 68704 561688 68710 561700
rect 69014 561688 69020 561700
rect 69072 561688 69078 561740
rect 4982 560260 4988 560312
rect 5040 560300 5046 560312
rect 67634 560300 67640 560312
rect 5040 560272 67640 560300
rect 5040 560260 5046 560272
rect 67634 560260 67640 560272
rect 67692 560260 67698 560312
rect 64874 559852 64880 559904
rect 64932 559892 64938 559904
rect 68646 559892 68652 559904
rect 64932 559864 68652 559892
rect 64932 559852 64938 559864
rect 68646 559852 68652 559864
rect 68704 559852 68710 559904
rect 57882 556180 57888 556232
rect 57940 556220 57946 556232
rect 64782 556220 64788 556232
rect 57940 556192 64788 556220
rect 57940 556180 57946 556192
rect 64782 556180 64788 556192
rect 64840 556180 64846 556232
rect 571334 554752 571340 554804
rect 571392 554792 571398 554804
rect 573726 554792 573732 554804
rect 571392 554764 573732 554792
rect 571392 554752 571398 554764
rect 573726 554752 573732 554764
rect 573784 554752 573790 554804
rect 55858 551760 55864 551812
rect 55916 551800 55922 551812
rect 57882 551800 57888 551812
rect 55916 551772 57888 551800
rect 55916 551760 55922 551772
rect 57882 551760 57888 551772
rect 57940 551760 57946 551812
rect 568942 548088 568948 548140
rect 569000 548128 569006 548140
rect 569402 548128 569408 548140
rect 569000 548100 569408 548128
rect 569000 548088 569006 548100
rect 569402 548088 569408 548100
rect 569460 548088 569466 548140
rect 55858 546496 55864 546508
rect 49712 546468 55864 546496
rect 47578 546388 47584 546440
rect 47636 546428 47642 546440
rect 49712 546428 49740 546468
rect 55858 546456 55864 546468
rect 55916 546456 55922 546508
rect 47636 546400 49740 546428
rect 47636 546388 47642 546400
rect 568942 540376 568948 540388
rect 568903 540348 568948 540376
rect 568942 540336 568948 540348
rect 569000 540336 569006 540388
rect 65978 536800 65984 536852
rect 66036 536840 66042 536852
rect 67634 536840 67640 536852
rect 66036 536812 67640 536840
rect 66036 536800 66042 536812
rect 67634 536800 67640 536812
rect 67692 536800 67698 536852
rect 42058 532040 42064 532092
rect 42116 532080 42122 532092
rect 47578 532080 47584 532092
rect 42116 532052 47584 532080
rect 42116 532040 42122 532052
rect 47578 532040 47584 532052
rect 47636 532040 47642 532092
rect 568942 525348 568948 525360
rect 568903 525320 568948 525348
rect 568942 525308 568948 525320
rect 569000 525308 569006 525360
rect 39666 514768 39672 514820
rect 39724 514808 39730 514820
rect 42058 514808 42064 514820
rect 39724 514780 42064 514808
rect 39724 514768 39730 514780
rect 42058 514768 42064 514780
rect 42116 514768 42122 514820
rect 571978 511912 571984 511964
rect 572036 511952 572042 511964
rect 580166 511952 580172 511964
rect 572036 511924 580172 511952
rect 572036 511912 572042 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 39666 510660 39672 510672
rect 37292 510632 39672 510660
rect 37182 510552 37188 510604
rect 37240 510592 37246 510604
rect 37292 510592 37320 510632
rect 39666 510620 39672 510632
rect 39724 510620 39730 510672
rect 37240 510564 37320 510592
rect 37240 510552 37246 510564
rect 568942 503044 568948 503056
rect 568903 503016 568948 503044
rect 568942 503004 568948 503016
rect 569000 503004 569006 503056
rect 35158 502936 35164 502988
rect 35216 502976 35222 502988
rect 37182 502976 37188 502988
rect 35216 502948 37188 502976
rect 35216 502936 35222 502948
rect 37182 502936 37188 502948
rect 37240 502936 37246 502988
rect 569034 499740 569040 499792
rect 569092 499780 569098 499792
rect 569402 499780 569408 499792
rect 569092 499752 569408 499780
rect 569092 499740 569098 499752
rect 569402 499740 569408 499752
rect 569460 499740 569466 499792
rect 568942 498080 568948 498092
rect 568868 498052 568948 498080
rect 568868 497808 568896 498052
rect 568942 498040 568948 498052
rect 569000 498040 569006 498092
rect 568942 497904 568948 497956
rect 569000 497944 569006 497956
rect 569402 497944 569408 497956
rect 569000 497916 569408 497944
rect 569000 497904 569006 497916
rect 569402 497904 569408 497916
rect 569460 497904 569466 497956
rect 568942 497808 568948 497820
rect 568868 497780 568948 497808
rect 568942 497768 568948 497780
rect 569000 497768 569006 497820
rect 568942 495360 568948 495372
rect 568903 495332 568948 495360
rect 568942 495320 568948 495332
rect 569000 495320 569006 495372
rect 33226 491240 33232 491292
rect 33284 491280 33290 491292
rect 35158 491280 35164 491292
rect 33284 491252 35164 491280
rect 33284 491240 33290 491252
rect 35158 491240 35164 491252
rect 35216 491240 35222 491292
rect 32398 487160 32404 487212
rect 32456 487200 32462 487212
rect 33226 487200 33232 487212
rect 32456 487172 33232 487200
rect 32456 487160 32462 487172
rect 33226 487160 33232 487172
rect 33284 487160 33290 487212
rect 568942 486452 568948 486464
rect 568903 486424 568948 486452
rect 568942 486412 568948 486424
rect 569000 486412 569006 486464
rect 568942 485092 568948 485104
rect 568903 485064 568948 485092
rect 568942 485052 568948 485064
rect 569000 485052 569006 485104
rect 30374 478864 30380 478916
rect 30432 478904 30438 478916
rect 32398 478904 32404 478916
rect 30432 478876 32404 478904
rect 30432 478864 30438 478876
rect 32398 478864 32404 478876
rect 32456 478864 32462 478916
rect 571334 477640 571340 477692
rect 571392 477680 571398 477692
rect 573634 477680 573640 477692
rect 571392 477652 573640 477680
rect 571392 477640 571398 477652
rect 573634 477640 573640 477652
rect 573692 477640 573698 477692
rect 2774 475872 2780 475924
rect 2832 475912 2838 475924
rect 5074 475912 5080 475924
rect 2832 475884 5080 475912
rect 2832 475872 2838 475884
rect 5074 475872 5080 475884
rect 5132 475872 5138 475924
rect 25130 469820 25136 469872
rect 25188 469860 25194 469872
rect 30006 469860 30012 469872
rect 25188 469832 30012 469860
rect 25188 469820 25194 469832
rect 30006 469820 30012 469832
rect 30064 469820 30070 469872
rect 24118 466420 24124 466472
rect 24176 466460 24182 466472
rect 25130 466460 25136 466472
rect 24176 466432 25136 466460
rect 24176 466420 24182 466432
rect 25130 466420 25136 466432
rect 25188 466420 25194 466472
rect 570598 458124 570604 458176
rect 570656 458164 570662 458176
rect 580166 458164 580172 458176
rect 570656 458136 580172 458164
rect 570656 458124 570662 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 68646 451120 68652 451172
rect 68704 451160 68710 451172
rect 69750 451160 69756 451172
rect 68704 451132 69756 451160
rect 68704 451120 68710 451132
rect 69750 451120 69756 451132
rect 69808 451120 69814 451172
rect 568942 445748 568948 445800
rect 569000 445788 569006 445800
rect 569402 445788 569408 445800
rect 569000 445760 569408 445788
rect 569000 445748 569006 445760
rect 569402 445748 569408 445760
rect 569460 445748 569466 445800
rect 568942 431536 568948 431588
rect 569000 431576 569006 431588
rect 569402 431576 569408 431588
rect 569000 431548 569408 431576
rect 569000 431536 569006 431548
rect 569402 431536 569408 431548
rect 569460 431536 569466 431588
rect 65794 426436 65800 426488
rect 65852 426476 65858 426488
rect 67910 426476 67916 426488
rect 65852 426448 67916 426476
rect 65852 426436 65858 426448
rect 67910 426436 67916 426448
rect 67968 426436 67974 426488
rect 22830 424736 22836 424788
rect 22888 424776 22894 424788
rect 24118 424776 24124 424788
rect 22888 424748 24124 424776
rect 22888 424736 22894 424748
rect 24118 424736 24124 424748
rect 24176 424736 24182 424788
rect 2774 423512 2780 423564
rect 2832 423552 2838 423564
rect 5074 423552 5080 423564
rect 2832 423524 5080 423552
rect 2832 423512 2838 423524
rect 5074 423512 5080 423524
rect 5132 423512 5138 423564
rect 575014 418140 575020 418192
rect 575072 418180 575078 418192
rect 580166 418180 580172 418192
rect 575072 418152 580172 418180
rect 575072 418140 575078 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 21358 417324 21364 417376
rect 21416 417364 21422 417376
rect 22830 417364 22836 417376
rect 21416 417336 22836 417364
rect 21416 417324 21422 417336
rect 22830 417324 22836 417336
rect 22888 417324 22894 417376
rect 13722 411272 13728 411324
rect 13780 411312 13786 411324
rect 67634 411312 67640 411324
rect 13780 411284 67640 411312
rect 13780 411272 13786 411284
rect 67634 411272 67640 411284
rect 67692 411272 67698 411324
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 50430 409884 50436 409896
rect 3384 409856 50436 409884
rect 3384 409844 3390 409856
rect 50430 409844 50436 409856
rect 50488 409844 50494 409896
rect 18598 408756 18604 408808
rect 18656 408796 18662 408808
rect 21358 408796 21364 408808
rect 18656 408768 21364 408796
rect 18656 408756 18662 408768
rect 21358 408756 21364 408768
rect 21416 408756 21422 408808
rect 15838 407192 15844 407244
rect 15896 407232 15902 407244
rect 18598 407232 18604 407244
rect 15896 407204 18604 407232
rect 15896 407192 15902 407204
rect 18598 407192 18604 407204
rect 18656 407192 18662 407244
rect 573726 405628 573732 405680
rect 573784 405668 573790 405680
rect 580166 405668 580172 405680
rect 573784 405640 580172 405668
rect 573784 405628 573790 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 65886 403248 65892 403300
rect 65944 403288 65950 403300
rect 68002 403288 68008 403300
rect 65944 403260 68008 403288
rect 65944 403248 65950 403260
rect 68002 403248 68008 403260
rect 68060 403248 68066 403300
rect 12434 400188 12440 400240
rect 12492 400228 12498 400240
rect 15838 400228 15844 400240
rect 12492 400200 15844 400228
rect 12492 400188 12498 400200
rect 15838 400188 15844 400200
rect 15896 400188 15902 400240
rect 5534 396720 5540 396772
rect 5592 396760 5598 396772
rect 12434 396760 12440 396772
rect 5592 396732 12440 396760
rect 5592 396720 5598 396732
rect 12434 396720 12440 396732
rect 12492 396720 12498 396772
rect 3970 396040 3976 396092
rect 4028 396080 4034 396092
rect 67634 396080 67640 396092
rect 4028 396052 67640 396080
rect 4028 396040 4034 396052
rect 67634 396040 67640 396052
rect 67692 396040 67698 396092
rect 569218 390532 569224 390584
rect 569276 390572 569282 390584
rect 571702 390572 571708 390584
rect 569276 390544 571708 390572
rect 569276 390532 569282 390544
rect 571702 390532 571708 390544
rect 571760 390532 571766 390584
rect 3694 372580 3700 372632
rect 3752 372620 3758 372632
rect 67634 372620 67640 372632
rect 3752 372592 67640 372620
rect 3752 372580 3758 372592
rect 67634 372580 67640 372592
rect 67692 372580 67698 372632
rect 3234 371220 3240 371272
rect 3292 371260 3298 371272
rect 5166 371260 5172 371272
rect 3292 371232 5172 371260
rect 3292 371220 3298 371232
rect 5166 371220 5172 371232
rect 5224 371220 5230 371272
rect 569310 365644 569316 365696
rect 569368 365684 569374 365696
rect 579982 365684 579988 365696
rect 569368 365656 579988 365684
rect 569368 365644 569374 365656
rect 579982 365644 579988 365656
rect 580040 365644 580046 365696
rect 55122 364352 55128 364404
rect 55180 364392 55186 364404
rect 67634 364392 67640 364404
rect 55180 364364 67640 364392
rect 55180 364352 55186 364364
rect 67634 364352 67640 364364
rect 67692 364352 67698 364404
rect 65702 356056 65708 356108
rect 65760 356096 65766 356108
rect 67818 356096 67824 356108
rect 65760 356068 67824 356096
rect 65760 356056 65766 356068
rect 67818 356056 67824 356068
rect 67876 356056 67882 356108
rect 3510 350480 3516 350532
rect 3568 350520 3574 350532
rect 67634 350520 67640 350532
rect 3568 350492 67640 350520
rect 3568 350480 3574 350492
rect 67634 350480 67640 350492
rect 67692 350480 67698 350532
rect 572070 344972 572076 345024
rect 572128 345012 572134 345024
rect 575014 345012 575020 345024
rect 572128 344984 575020 345012
rect 572128 344972 572134 344984
rect 575014 344972 575020 344984
rect 575072 344972 575078 345024
rect 52362 342864 52368 342916
rect 52420 342904 52426 342916
rect 65518 342904 65524 342916
rect 52420 342876 65524 342904
rect 52420 342864 52426 342876
rect 65518 342864 65524 342876
rect 65576 342864 65582 342916
rect 572622 329536 572628 329588
rect 572680 329576 572686 329588
rect 576210 329576 576216 329588
rect 572680 329548 576216 329576
rect 572680 329536 572686 329548
rect 576210 329536 576216 329548
rect 576268 329536 576274 329588
rect 24762 327020 24768 327072
rect 24820 327060 24826 327072
rect 67634 327060 67640 327072
rect 24820 327032 67640 327060
rect 24820 327020 24826 327032
rect 67634 327020 67640 327032
rect 67692 327020 67698 327072
rect 568942 321580 568948 321632
rect 569000 321620 569006 321632
rect 569310 321620 569316 321632
rect 569000 321592 569316 321620
rect 569000 321580 569006 321592
rect 569310 321580 569316 321592
rect 569368 321580 569374 321632
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 7650 320124 7656 320136
rect 3568 320096 7656 320124
rect 3568 320084 3574 320096
rect 7650 320084 7656 320096
rect 7708 320084 7714 320136
rect 68186 310428 68192 310480
rect 68244 310468 68250 310480
rect 69842 310468 69848 310480
rect 68244 310440 69848 310468
rect 68244 310428 68250 310440
rect 69842 310428 69848 310440
rect 69900 310428 69906 310480
rect 571334 305600 571340 305652
rect 571392 305640 571398 305652
rect 572990 305640 572996 305652
rect 571392 305612 572996 305640
rect 571392 305600 571398 305612
rect 572990 305600 572996 305612
rect 573048 305600 573054 305652
rect 27522 302880 27528 302932
rect 27580 302920 27586 302932
rect 68278 302920 68284 302932
rect 27580 302892 68284 302920
rect 27580 302880 27586 302892
rect 68278 302880 68284 302892
rect 68336 302880 68342 302932
rect 65518 302200 65524 302252
rect 65576 302240 65582 302252
rect 67818 302240 67824 302252
rect 65576 302212 67824 302240
rect 65576 302200 65582 302212
rect 67818 302200 67824 302212
rect 67876 302200 67882 302252
rect 576302 299412 576308 299464
rect 576360 299452 576366 299464
rect 580166 299452 580172 299464
rect 576360 299424 580172 299452
rect 576360 299412 576366 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 65610 285676 65616 285728
rect 65668 285716 65674 285728
rect 67818 285716 67824 285728
rect 65668 285688 67824 285716
rect 65668 285676 65674 285688
rect 67818 285676 67824 285688
rect 67876 285676 67882 285728
rect 3878 270512 3884 270564
rect 3936 270552 3942 270564
rect 67634 270552 67640 270564
rect 3936 270524 67640 270552
rect 3936 270512 3942 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 569034 266364 569040 266416
rect 569092 266404 569098 266416
rect 569310 266404 569316 266416
rect 569092 266376 569316 266404
rect 569092 266364 569098 266376
rect 569310 266364 569316 266376
rect 569368 266364 569374 266416
rect 569126 258476 569132 258528
rect 569184 258516 569190 258528
rect 569310 258516 569316 258528
rect 569184 258488 569316 258516
rect 569184 258476 569190 258488
rect 569310 258476 569316 258488
rect 569368 258476 569374 258528
rect 575014 258068 575020 258120
rect 575072 258108 575078 258120
rect 579614 258108 579620 258120
rect 575072 258080 579620 258108
rect 575072 258068 575078 258080
rect 579614 258068 579620 258080
rect 579672 258068 579678 258120
rect 68370 247664 68376 247716
rect 68428 247704 68434 247716
rect 69842 247704 69848 247716
rect 68428 247676 69848 247704
rect 68428 247664 68434 247676
rect 69842 247664 69848 247676
rect 69900 247664 69906 247716
rect 574922 245556 574928 245608
rect 574980 245596 574986 245608
rect 580166 245596 580172 245608
rect 574980 245568 580172 245596
rect 574980 245556 574986 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 63402 238756 63408 238808
rect 63460 238796 63466 238808
rect 67634 238796 67640 238808
rect 63460 238768 67640 238796
rect 63460 238756 63466 238768
rect 67634 238756 67640 238768
rect 67692 238756 67698 238808
rect 10962 231820 10968 231872
rect 11020 231860 11026 231872
rect 67634 231860 67640 231872
rect 11020 231832 67640 231860
rect 11020 231820 11026 231832
rect 67634 231820 67640 231832
rect 67692 231820 67698 231872
rect 568942 219716 568948 219768
rect 569000 219756 569006 219768
rect 569402 219756 569408 219768
rect 569000 219728 569408 219756
rect 569000 219716 569006 219728
rect 569402 219716 569408 219728
rect 569460 219716 569466 219768
rect 574922 218016 574928 218068
rect 574980 218056 574986 218068
rect 580166 218056 580172 218068
rect 574980 218028 580172 218056
rect 574980 218016 574986 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 26142 208360 26148 208412
rect 26200 208400 26206 208412
rect 67634 208400 67640 208412
rect 26200 208372 67640 208400
rect 26200 208360 26206 208372
rect 67634 208360 67640 208372
rect 67692 208360 67698 208412
rect 68370 193128 68376 193180
rect 68428 193168 68434 193180
rect 69566 193168 69572 193180
rect 68428 193140 69572 193168
rect 68428 193128 68434 193140
rect 69566 193128 69572 193140
rect 69624 193128 69630 193180
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 5166 187728 5172 187740
rect 3384 187700 5172 187728
rect 3384 187688 3390 187700
rect 5166 187688 5172 187700
rect 5224 187688 5230 187740
rect 577498 179324 577504 179376
rect 577556 179364 577562 179376
rect 579890 179364 579896 179376
rect 577556 179336 579896 179364
rect 577556 179324 577562 179336
rect 579890 179324 579896 179336
rect 579948 179324 579954 179376
rect 9582 176672 9588 176724
rect 9640 176712 9646 176724
rect 67634 176712 67640 176724
rect 9640 176684 67640 176712
rect 9640 176672 9646 176684
rect 67634 176672 67640 176684
rect 67692 176672 67698 176724
rect 5534 171096 5540 171148
rect 5592 171136 5598 171148
rect 5592 171108 6960 171136
rect 5592 171096 5598 171108
rect 6932 171068 6960 171108
rect 8294 171068 8300 171080
rect 6932 171040 8300 171068
rect 8294 171028 8300 171040
rect 8352 171028 8358 171080
rect 8294 168376 8300 168428
rect 8352 168416 8358 168428
rect 9766 168416 9772 168428
rect 8352 168388 9772 168416
rect 8352 168376 8358 168388
rect 9766 168376 9772 168388
rect 9824 168376 9830 168428
rect 574830 166948 574836 167000
rect 574888 166988 574894 167000
rect 580166 166988 580172 167000
rect 574888 166960 580172 166988
rect 574888 166948 574894 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 9766 164228 9772 164280
rect 9824 164268 9830 164280
rect 9824 164240 11100 164268
rect 9824 164228 9830 164240
rect 11072 164200 11100 164240
rect 15194 164200 15200 164212
rect 11072 164172 15200 164200
rect 15194 164160 15200 164172
rect 15252 164160 15258 164212
rect 65426 161508 65432 161560
rect 65484 161548 65490 161560
rect 67634 161548 67640 161560
rect 65484 161520 67640 161548
rect 65484 161508 65490 161520
rect 67634 161508 67640 161520
rect 67692 161508 67698 161560
rect 15194 161372 15200 161424
rect 15252 161412 15258 161424
rect 19242 161412 19248 161424
rect 15252 161384 19248 161412
rect 15252 161372 15258 161384
rect 19242 161372 19248 161384
rect 19300 161372 19306 161424
rect 19334 151784 19340 151836
rect 19392 151824 19398 151836
rect 19392 151796 20760 151824
rect 19392 151784 19398 151796
rect 20732 151756 20760 151796
rect 22830 151756 22836 151768
rect 20732 151728 22836 151756
rect 22830 151716 22836 151728
rect 22888 151716 22894 151768
rect 2774 150084 2780 150136
rect 2832 150124 2838 150136
rect 4982 150124 4988 150136
rect 2832 150096 4988 150124
rect 2832 150084 2838 150096
rect 4982 150084 4988 150096
rect 5040 150084 5046 150136
rect 68094 146208 68100 146260
rect 68152 146248 68158 146260
rect 69474 146248 69480 146260
rect 68152 146220 69480 146248
rect 68152 146208 68158 146220
rect 69474 146208 69480 146220
rect 69532 146208 69538 146260
rect 570782 140768 570788 140820
rect 570840 140808 570846 140820
rect 571794 140808 571800 140820
rect 570840 140780 571800 140808
rect 570840 140768 570846 140780
rect 571794 140768 571800 140780
rect 571852 140768 571858 140820
rect 3602 139340 3608 139392
rect 3660 139380 3666 139392
rect 67634 139380 67640 139392
rect 3660 139352 67640 139380
rect 3660 139340 3666 139352
rect 67634 139340 67640 139352
rect 67692 139340 67698 139392
rect 573634 139340 573640 139392
rect 573692 139380 573698 139392
rect 580166 139380 580172 139392
rect 573692 139352 580172 139380
rect 573692 139340 573698 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 22830 138660 22836 138712
rect 22888 138700 22894 138712
rect 24118 138700 24124 138712
rect 22888 138672 24124 138700
rect 22888 138660 22894 138672
rect 24118 138660 24124 138672
rect 24176 138660 24182 138712
rect 24118 129752 24124 129804
rect 24176 129792 24182 129804
rect 24176 129764 26234 129792
rect 24176 129752 24182 129764
rect 26206 129724 26234 129764
rect 66806 129752 66812 129804
rect 66864 129792 66870 129804
rect 67634 129792 67640 129804
rect 66864 129764 67640 129792
rect 66864 129752 66870 129764
rect 67634 129752 67640 129764
rect 67692 129752 67698 129804
rect 28258 129724 28264 129736
rect 26206 129696 28264 129724
rect 28258 129684 28264 129696
rect 28316 129684 28322 129736
rect 573542 126896 573548 126948
rect 573600 126936 573606 126948
rect 579614 126936 579620 126948
rect 573600 126908 579620 126936
rect 573600 126896 573606 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 28258 125536 28264 125588
rect 28316 125576 28322 125588
rect 30282 125576 30288 125588
rect 28316 125548 30288 125576
rect 28316 125536 28322 125548
rect 30282 125536 30288 125548
rect 30340 125536 30346 125588
rect 30374 118124 30380 118176
rect 30432 118164 30438 118176
rect 32398 118164 32404 118176
rect 30432 118136 32404 118164
rect 30432 118124 30438 118136
rect 32398 118124 32404 118136
rect 32456 118124 32462 118176
rect 32398 105476 32404 105528
rect 32456 105516 32462 105528
rect 37274 105516 37280 105528
rect 32456 105488 37280 105516
rect 32456 105476 32462 105488
rect 37274 105476 37280 105488
rect 37332 105476 37338 105528
rect 37274 100852 37280 100904
rect 37332 100892 37338 100904
rect 40034 100892 40040 100904
rect 37332 100864 40040 100892
rect 37332 100852 37338 100864
rect 40034 100852 40040 100864
rect 40092 100852 40098 100904
rect 576118 100648 576124 100700
rect 576176 100688 576182 100700
rect 579706 100688 579712 100700
rect 576176 100660 579712 100688
rect 576176 100648 576182 100660
rect 579706 100648 579712 100660
rect 579764 100648 579770 100700
rect 22002 97996 22008 98048
rect 22060 98036 22066 98048
rect 67634 98036 67640 98048
rect 22060 98008 67640 98036
rect 22060 97996 22066 98008
rect 67634 97996 67640 98008
rect 67692 97996 67698 98048
rect 3326 97928 3332 97980
rect 3384 97968 3390 97980
rect 10410 97968 10416 97980
rect 3384 97940 10416 97968
rect 3384 97928 3390 97940
rect 10410 97928 10416 97940
rect 10468 97928 10474 97980
rect 40034 95140 40040 95192
rect 40092 95180 40098 95192
rect 42610 95180 42616 95192
rect 40092 95152 42616 95180
rect 40092 95140 40098 95152
rect 42610 95140 42616 95152
rect 42668 95140 42674 95192
rect 42610 92284 42616 92336
rect 42668 92324 42674 92336
rect 44174 92324 44180 92336
rect 42668 92296 44180 92324
rect 42668 92284 42674 92296
rect 44174 92284 44180 92296
rect 44232 92284 44238 92336
rect 44174 90312 44180 90364
rect 44232 90352 44238 90364
rect 49602 90352 49608 90364
rect 44232 90324 49608 90352
rect 44232 90312 44238 90324
rect 49602 90312 49608 90324
rect 49660 90312 49666 90364
rect 49694 86912 49700 86964
rect 49752 86952 49758 86964
rect 52270 86952 52276 86964
rect 49752 86924 52276 86952
rect 49752 86912 49758 86924
rect 52270 86912 52276 86924
rect 52328 86912 52334 86964
rect 37182 82832 37188 82884
rect 37240 82872 37246 82884
rect 68370 82872 68376 82884
rect 37240 82844 68376 82872
rect 37240 82832 37246 82844
rect 68370 82832 68376 82844
rect 68428 82832 68434 82884
rect 52270 82424 52276 82476
rect 52328 82464 52334 82476
rect 56502 82464 56508 82476
rect 52328 82436 56508 82464
rect 52328 82424 52334 82436
rect 56502 82424 56508 82436
rect 56560 82424 56566 82476
rect 569770 80044 569776 80096
rect 569828 80084 569834 80096
rect 571518 80084 571524 80096
rect 569828 80056 571524 80084
rect 569828 80044 569834 80056
rect 571518 80044 571524 80056
rect 571576 80044 571582 80096
rect 56502 77256 56508 77308
rect 56560 77296 56566 77308
rect 56560 77268 58020 77296
rect 56560 77256 56566 77268
rect 57992 77228 58020 77268
rect 63494 77228 63500 77240
rect 57992 77200 63500 77228
rect 63494 77188 63500 77200
rect 63552 77188 63558 77240
rect 63494 75148 63500 75200
rect 63552 75188 63558 75200
rect 69382 75188 69388 75200
rect 63552 75160 69388 75188
rect 63552 75148 63558 75160
rect 69382 75148 69388 75160
rect 69440 75148 69446 75200
rect 569310 71136 569316 71188
rect 569368 71176 569374 71188
rect 569862 71176 569868 71188
rect 569368 71148 569868 71176
rect 569368 71136 569374 71148
rect 569862 71136 569868 71148
rect 569920 71136 569926 71188
rect 50982 70048 50988 70100
rect 51040 70088 51046 70100
rect 570598 70088 570604 70100
rect 51040 70060 570604 70088
rect 51040 70048 51046 70060
rect 570598 70048 570604 70060
rect 570656 70048 570662 70100
rect 42702 69980 42708 70032
rect 42760 70020 42766 70032
rect 570322 70020 570328 70032
rect 42760 69992 570328 70020
rect 42760 69980 42766 69992
rect 570322 69980 570328 69992
rect 570380 69980 570386 70032
rect 37090 69912 37096 69964
rect 37148 69952 37154 69964
rect 570506 69952 570512 69964
rect 37148 69924 570512 69952
rect 37148 69912 37154 69924
rect 570506 69912 570512 69924
rect 570564 69912 570570 69964
rect 35802 69844 35808 69896
rect 35860 69884 35866 69896
rect 570966 69884 570972 69896
rect 35860 69856 570972 69884
rect 35860 69844 35866 69856
rect 570966 69844 570972 69856
rect 571024 69844 571030 69896
rect 21358 69776 21364 69828
rect 21416 69816 21422 69828
rect 567749 69819 567807 69825
rect 567749 69816 567761 69819
rect 21416 69788 567761 69816
rect 21416 69776 21422 69788
rect 567749 69785 567761 69788
rect 567795 69785 567807 69819
rect 567749 69779 567807 69785
rect 567838 69776 567844 69828
rect 567896 69816 567902 69828
rect 571978 69816 571984 69828
rect 567896 69788 571984 69816
rect 567896 69776 567902 69788
rect 571978 69776 571984 69788
rect 572036 69776 572042 69828
rect 7650 69708 7656 69760
rect 7708 69748 7714 69760
rect 572070 69748 572076 69760
rect 7708 69720 572076 69748
rect 7708 69708 7714 69720
rect 572070 69708 572076 69720
rect 572128 69708 572134 69760
rect 4982 69640 4988 69692
rect 5040 69680 5046 69692
rect 571334 69680 571340 69692
rect 5040 69652 571340 69680
rect 5040 69640 5046 69652
rect 571334 69640 571340 69652
rect 571392 69640 571398 69692
rect 57882 69572 57888 69624
rect 57940 69612 57946 69624
rect 571426 69612 571432 69624
rect 57940 69584 571432 69612
rect 57940 69572 57946 69584
rect 571426 69572 571432 69584
rect 571484 69572 571490 69624
rect 69014 69504 69020 69556
rect 69072 69544 69078 69556
rect 580534 69544 580540 69556
rect 69072 69516 580540 69544
rect 69072 69504 69078 69516
rect 580534 69504 580540 69516
rect 580592 69504 580598 69556
rect 67634 69436 67640 69488
rect 67692 69476 67698 69488
rect 580258 69476 580264 69488
rect 67692 69448 580264 69476
rect 67692 69436 67698 69448
rect 580258 69436 580264 69448
rect 580316 69436 580322 69488
rect 61930 69368 61936 69420
rect 61988 69408 61994 69420
rect 567657 69411 567715 69417
rect 567657 69408 567669 69411
rect 61988 69380 567669 69408
rect 61988 69368 61994 69380
rect 567657 69377 567669 69380
rect 567703 69377 567715 69411
rect 567657 69371 567715 69377
rect 567749 69411 567807 69417
rect 567749 69377 567761 69411
rect 567795 69408 567807 69411
rect 572254 69408 572260 69420
rect 567795 69380 572260 69408
rect 567795 69377 567807 69380
rect 567749 69371 567807 69377
rect 572254 69368 572260 69380
rect 572312 69368 572318 69420
rect 65334 69300 65340 69352
rect 65392 69340 65398 69352
rect 569034 69340 569040 69352
rect 65392 69312 569040 69340
rect 65392 69300 65398 69312
rect 569034 69300 569040 69312
rect 569092 69300 569098 69352
rect 69382 69232 69388 69284
rect 69440 69272 69446 69284
rect 569586 69272 569592 69284
rect 69440 69244 569592 69272
rect 69440 69232 69446 69244
rect 569586 69232 569592 69244
rect 569644 69232 569650 69284
rect 567657 69207 567715 69213
rect 567657 69173 567669 69207
rect 567703 69204 567715 69207
rect 571886 69204 571892 69216
rect 567703 69176 571892 69204
rect 567703 69173 567715 69176
rect 567657 69167 567715 69173
rect 571886 69164 571892 69176
rect 571944 69164 571950 69216
rect 68738 69136 68744 69148
rect 68664 69108 68744 69136
rect 68370 68960 68376 69012
rect 68428 69000 68434 69012
rect 68664 69000 68692 69108
rect 68738 69096 68744 69108
rect 68796 69096 68802 69148
rect 68428 68972 68692 69000
rect 68428 68960 68434 68972
rect 68738 68960 68744 69012
rect 68796 69000 68802 69012
rect 68922 69000 68928 69012
rect 68796 68972 68928 69000
rect 68796 68960 68802 68972
rect 68922 68960 68928 68972
rect 68980 68960 68986 69012
rect 69017 69003 69075 69009
rect 69017 68969 69029 69003
rect 69063 69000 69075 69003
rect 197357 69003 197415 69009
rect 197357 69000 197369 69003
rect 69063 68972 197369 69000
rect 69063 68969 69075 68972
rect 69017 68963 69075 68969
rect 197357 68969 197369 68972
rect 197403 68969 197415 69003
rect 197357 68963 197415 68969
rect 200025 69003 200083 69009
rect 200025 68969 200037 69003
rect 200071 69000 200083 69003
rect 569402 69000 569408 69012
rect 200071 68972 569408 69000
rect 200071 68969 200083 68972
rect 200025 68963 200083 68969
rect 569402 68960 569408 68972
rect 569460 68960 569466 69012
rect 67726 68892 67732 68944
rect 67784 68932 67790 68944
rect 178037 68935 178095 68941
rect 178037 68932 178049 68935
rect 67784 68904 178049 68932
rect 67784 68892 67790 68904
rect 178037 68901 178049 68904
rect 178083 68901 178095 68935
rect 178037 68895 178095 68901
rect 190365 68935 190423 68941
rect 190365 68901 190377 68935
rect 190411 68932 190423 68935
rect 570414 68932 570420 68944
rect 190411 68904 570420 68932
rect 190411 68901 190423 68904
rect 190365 68895 190423 68901
rect 570414 68892 570420 68904
rect 570472 68892 570478 68944
rect 67910 68824 67916 68876
rect 67968 68864 67974 68876
rect 182177 68867 182235 68873
rect 182177 68864 182189 68867
rect 67968 68836 182189 68864
rect 67968 68824 67974 68836
rect 182177 68833 182189 68836
rect 182223 68833 182235 68867
rect 182177 68827 182235 68833
rect 186041 68867 186099 68873
rect 186041 68833 186053 68867
rect 186087 68864 186099 68867
rect 569678 68864 569684 68876
rect 186087 68836 569684 68864
rect 186087 68833 186099 68836
rect 186041 68827 186099 68833
rect 569678 68824 569684 68836
rect 569736 68824 569742 68876
rect 68922 68756 68928 68808
rect 68980 68796 68986 68808
rect 69658 68796 69664 68808
rect 68980 68768 69664 68796
rect 68980 68756 68986 68768
rect 69658 68756 69664 68768
rect 69716 68756 69722 68808
rect 154301 68799 154359 68805
rect 154301 68765 154313 68799
rect 154347 68796 154359 68799
rect 569954 68796 569960 68808
rect 154347 68768 569960 68796
rect 154347 68765 154359 68768
rect 154301 68759 154359 68765
rect 569954 68756 569960 68768
rect 570012 68756 570018 68808
rect 66990 68688 66996 68740
rect 67048 68728 67054 68740
rect 69017 68731 69075 68737
rect 69017 68728 69029 68731
rect 67048 68700 69029 68728
rect 67048 68688 67054 68700
rect 69017 68697 69029 68700
rect 69063 68697 69075 68731
rect 69017 68691 69075 68697
rect 69290 68688 69296 68740
rect 69348 68728 69354 68740
rect 70394 68728 70400 68740
rect 69348 68700 70400 68728
rect 69348 68688 69354 68700
rect 70394 68688 70400 68700
rect 70452 68688 70458 68740
rect 132586 68728 132592 68740
rect 70596 68700 132592 68728
rect 68554 68620 68560 68672
rect 68612 68660 68618 68672
rect 70596 68660 70624 68700
rect 132586 68688 132592 68700
rect 132644 68688 132650 68740
rect 153102 68688 153108 68740
rect 153160 68728 153166 68740
rect 572530 68728 572536 68740
rect 153160 68700 572536 68728
rect 153160 68688 153166 68700
rect 572530 68688 572536 68700
rect 572588 68688 572594 68740
rect 140774 68660 140780 68672
rect 68612 68632 70624 68660
rect 72528 68632 140780 68660
rect 68612 68620 68618 68632
rect 67818 68552 67824 68604
rect 67876 68592 67882 68604
rect 72418 68592 72424 68604
rect 67876 68564 72424 68592
rect 67876 68552 67882 68564
rect 72418 68552 72424 68564
rect 72476 68552 72482 68604
rect 66806 68484 66812 68536
rect 66864 68524 66870 68536
rect 72528 68524 72556 68632
rect 140774 68620 140780 68632
rect 140832 68620 140838 68672
rect 152093 68663 152151 68669
rect 152093 68629 152105 68663
rect 152139 68660 152151 68663
rect 572438 68660 572444 68672
rect 152139 68632 572444 68660
rect 152139 68629 152151 68632
rect 152093 68623 152151 68629
rect 572438 68620 572444 68632
rect 572496 68620 572502 68672
rect 128354 68552 128360 68604
rect 128412 68592 128418 68604
rect 570230 68592 570236 68604
rect 128412 68564 570236 68592
rect 128412 68552 128418 68564
rect 570230 68552 570236 68564
rect 570288 68552 570294 68604
rect 66864 68496 72556 68524
rect 72605 68527 72663 68533
rect 66864 68484 66870 68496
rect 72605 68493 72617 68527
rect 72651 68524 72663 68527
rect 84194 68524 84200 68536
rect 72651 68496 84200 68524
rect 72651 68493 72663 68496
rect 72605 68487 72663 68493
rect 84194 68484 84200 68496
rect 84252 68484 84258 68536
rect 126882 68484 126888 68536
rect 126940 68524 126946 68536
rect 570046 68524 570052 68536
rect 126940 68496 570052 68524
rect 126940 68484 126946 68496
rect 570046 68484 570052 68496
rect 570104 68484 570110 68536
rect 68830 68416 68836 68468
rect 68888 68456 68894 68468
rect 80146 68456 80152 68468
rect 68888 68428 80152 68456
rect 68888 68416 68894 68428
rect 80146 68416 80152 68428
rect 80204 68416 80210 68468
rect 84102 68416 84108 68468
rect 84160 68456 84166 68468
rect 568666 68456 568672 68468
rect 84160 68428 568672 68456
rect 84160 68416 84166 68428
rect 568666 68416 568672 68428
rect 568724 68416 568730 68468
rect 66070 68348 66076 68400
rect 66128 68388 66134 68400
rect 73154 68388 73160 68400
rect 66128 68360 73160 68388
rect 66128 68348 66134 68360
rect 73154 68348 73160 68360
rect 73212 68348 73218 68400
rect 77202 68348 77208 68400
rect 77260 68388 77266 68400
rect 569310 68388 569316 68400
rect 77260 68360 569316 68388
rect 77260 68348 77266 68360
rect 569310 68348 569316 68360
rect 569368 68348 569374 68400
rect 65702 68280 65708 68332
rect 65760 68320 65766 68332
rect 72605 68323 72663 68329
rect 72605 68320 72617 68323
rect 65760 68292 72617 68320
rect 65760 68280 65766 68292
rect 72605 68289 72617 68292
rect 72651 68289 72663 68323
rect 72605 68283 72663 68289
rect 73062 68280 73068 68332
rect 73120 68320 73126 68332
rect 572162 68320 572168 68332
rect 73120 68292 572168 68320
rect 73120 68280 73126 68292
rect 572162 68280 572168 68292
rect 572220 68280 572226 68332
rect 66898 68212 66904 68264
rect 66956 68252 66962 68264
rect 190546 68252 190552 68264
rect 66956 68224 190552 68252
rect 66956 68212 66962 68224
rect 190546 68212 190552 68224
rect 190604 68212 190610 68264
rect 197354 68252 197360 68264
rect 197315 68224 197360 68252
rect 197354 68212 197360 68224
rect 197412 68212 197418 68264
rect 200022 68252 200028 68264
rect 199983 68224 200028 68252
rect 200022 68212 200028 68224
rect 200080 68212 200086 68264
rect 206922 68212 206928 68264
rect 206980 68252 206986 68264
rect 571794 68252 571800 68264
rect 206980 68224 571800 68252
rect 206980 68212 206986 68224
rect 571794 68212 571800 68224
rect 571852 68212 571858 68264
rect 67174 68144 67180 68196
rect 67232 68184 67238 68196
rect 211154 68184 211160 68196
rect 67232 68156 211160 68184
rect 67232 68144 67238 68156
rect 211154 68144 211160 68156
rect 211212 68144 211218 68196
rect 219342 68144 219348 68196
rect 219400 68184 219406 68196
rect 570690 68184 570696 68196
rect 219400 68156 570696 68184
rect 219400 68144 219406 68156
rect 570690 68144 570696 68156
rect 570748 68144 570754 68196
rect 67358 68076 67364 68128
rect 67416 68116 67422 68128
rect 222194 68116 222200 68128
rect 67416 68088 222200 68116
rect 67416 68076 67422 68088
rect 222194 68076 222200 68088
rect 222252 68076 222258 68128
rect 226242 68076 226248 68128
rect 226300 68116 226306 68128
rect 570138 68116 570144 68128
rect 226300 68088 570144 68116
rect 226300 68076 226306 68088
rect 570138 68076 570144 68088
rect 570196 68076 570202 68128
rect 68738 68008 68744 68060
rect 68796 68048 68802 68060
rect 227806 68048 227812 68060
rect 68796 68020 227812 68048
rect 68796 68008 68802 68020
rect 227806 68008 227812 68020
rect 227864 68008 227870 68060
rect 230382 68008 230388 68060
rect 230440 68048 230446 68060
rect 569126 68048 569132 68060
rect 230440 68020 569132 68048
rect 230440 68008 230446 68020
rect 569126 68008 569132 68020
rect 569184 68008 569190 68060
rect 69198 67940 69204 67992
rect 69256 67980 69262 67992
rect 74626 67980 74632 67992
rect 69256 67952 74632 67980
rect 69256 67940 69262 67952
rect 74626 67940 74632 67952
rect 74684 67940 74690 67992
rect 79321 67983 79379 67989
rect 79321 67949 79333 67983
rect 79367 67980 79379 67983
rect 220814 67980 220820 67992
rect 79367 67952 220820 67980
rect 79367 67949 79379 67952
rect 79321 67943 79379 67949
rect 220814 67940 220820 67952
rect 220872 67940 220878 67992
rect 65794 67872 65800 67924
rect 65852 67912 65858 67924
rect 209774 67912 209780 67924
rect 65852 67884 209780 67912
rect 65852 67872 65858 67884
rect 209774 67872 209780 67884
rect 209832 67872 209838 67924
rect 65426 67804 65432 67856
rect 65484 67844 65490 67856
rect 166994 67844 167000 67856
rect 65484 67816 167000 67844
rect 65484 67804 65490 67816
rect 166994 67804 167000 67816
rect 167052 67804 167058 67856
rect 178034 67844 178040 67856
rect 177995 67816 178040 67844
rect 178034 67804 178040 67816
rect 178092 67804 178098 67856
rect 182174 67844 182180 67856
rect 182135 67816 182180 67844
rect 182174 67804 182180 67816
rect 182232 67804 182238 67856
rect 186038 67844 186044 67856
rect 185999 67816 186044 67844
rect 186038 67804 186044 67816
rect 186096 67804 186102 67856
rect 190362 67844 190368 67856
rect 190323 67816 190368 67844
rect 190362 67804 190368 67816
rect 190420 67804 190426 67856
rect 67266 67736 67272 67788
rect 67324 67776 67330 67788
rect 161474 67776 161480 67788
rect 67324 67748 161480 67776
rect 67324 67736 67330 67748
rect 161474 67736 161480 67748
rect 161532 67736 161538 67788
rect 68002 67668 68008 67720
rect 68060 67708 68066 67720
rect 157334 67708 157340 67720
rect 68060 67680 157340 67708
rect 68060 67668 68066 67680
rect 157334 67668 157340 67680
rect 157392 67668 157398 67720
rect 68370 67600 68376 67652
rect 68428 67640 68434 67652
rect 79321 67643 79379 67649
rect 79321 67640 79333 67643
rect 68428 67612 79333 67640
rect 68428 67600 68434 67612
rect 79321 67609 79333 67612
rect 79367 67609 79379 67643
rect 79321 67603 79379 67609
rect 150342 67600 150348 67652
rect 150400 67640 150406 67652
rect 152093 67643 152151 67649
rect 152093 67640 152105 67643
rect 150400 67612 152105 67640
rect 150400 67600 150406 67612
rect 152093 67609 152105 67612
rect 152139 67609 152151 67643
rect 154298 67640 154304 67652
rect 154259 67612 154304 67640
rect 152093 67603 152151 67609
rect 154298 67600 154304 67612
rect 154356 67600 154362 67652
rect 4890 67532 4896 67584
rect 4948 67572 4954 67584
rect 545850 67572 545856 67584
rect 4948 67544 545856 67572
rect 4948 67532 4954 67544
rect 545850 67532 545856 67544
rect 545908 67532 545914 67584
rect 4798 67464 4804 67516
rect 4856 67504 4862 67516
rect 503530 67504 503536 67516
rect 4856 67476 503536 67504
rect 4856 67464 4862 67476
rect 503530 67464 503536 67476
rect 503588 67464 503594 67516
rect 4062 67396 4068 67448
rect 4120 67436 4126 67448
rect 477034 67436 477040 67448
rect 4120 67408 477040 67436
rect 4120 67396 4126 67408
rect 477034 67396 477040 67408
rect 477092 67396 477098 67448
rect 7558 67328 7564 67380
rect 7616 67368 7622 67380
rect 418890 67368 418896 67380
rect 7616 67340 418896 67368
rect 7616 67328 7622 67340
rect 418890 67328 418896 67340
rect 418948 67328 418954 67380
rect 3786 67260 3792 67312
rect 3844 67300 3850 67312
rect 387242 67300 387248 67312
rect 3844 67272 387248 67300
rect 3844 67260 3850 67272
rect 387242 67260 387248 67272
rect 387300 67260 387306 67312
rect 5074 67192 5080 67244
rect 5132 67232 5138 67244
rect 128170 67232 128176 67244
rect 5132 67204 128176 67232
rect 5132 67192 5138 67204
rect 128170 67192 128176 67204
rect 128228 67192 128234 67244
rect 366082 67192 366088 67244
rect 366140 67232 366146 67244
rect 574922 67232 574928 67244
rect 366140 67204 574928 67232
rect 366140 67192 366146 67204
rect 574922 67192 574928 67204
rect 574980 67192 574986 67244
rect 119982 67124 119988 67176
rect 120040 67164 120046 67176
rect 572346 67164 572352 67176
rect 120040 67136 572352 67164
rect 120040 67124 120046 67136
rect 572346 67124 572352 67136
rect 572404 67124 572410 67176
rect 115842 67056 115848 67108
rect 115900 67096 115906 67108
rect 568758 67096 568764 67108
rect 115900 67068 568764 67096
rect 115900 67056 115906 67068
rect 568758 67056 568764 67068
rect 568816 67056 568822 67108
rect 65978 66988 65984 67040
rect 66036 67028 66042 67040
rect 91094 67028 91100 67040
rect 66036 67000 91100 67028
rect 66036 66988 66042 67000
rect 91094 66988 91100 67000
rect 91152 66988 91158 67040
rect 111702 66988 111708 67040
rect 111760 67028 111766 67040
rect 569862 67028 569868 67040
rect 111760 67000 569868 67028
rect 111760 66988 111766 67000
rect 569862 66988 569868 67000
rect 569920 66988 569926 67040
rect 67082 66920 67088 66972
rect 67140 66960 67146 66972
rect 580258 66960 580264 66972
rect 67140 66932 580264 66960
rect 67140 66920 67146 66932
rect 580258 66920 580264 66932
rect 580316 66920 580322 66972
rect 3694 66852 3700 66904
rect 3752 66892 3758 66904
rect 570874 66892 570880 66904
rect 3752 66864 570880 66892
rect 3752 66852 3758 66864
rect 570874 66852 570880 66864
rect 570932 66852 570938 66904
rect 3510 66784 3516 66836
rect 3568 66824 3574 66836
rect 175642 66824 175648 66836
rect 3568 66796 175648 66824
rect 3568 66784 3574 66796
rect 175642 66784 175648 66796
rect 175700 66784 175706 66836
rect 254946 66784 254952 66836
rect 255004 66824 255010 66836
rect 580350 66824 580356 66836
rect 255004 66796 580356 66824
rect 255004 66784 255010 66796
rect 580350 66784 580356 66796
rect 580408 66784 580414 66836
rect 67450 66716 67456 66768
rect 67508 66756 67514 66768
rect 208394 66756 208400 66768
rect 67508 66728 208400 66756
rect 67508 66716 67514 66728
rect 208394 66716 208400 66728
rect 208452 66716 208458 66768
rect 260282 66716 260288 66768
rect 260340 66756 260346 66768
rect 580442 66756 580448 66768
rect 260340 66728 580448 66756
rect 260340 66716 260346 66728
rect 580442 66716 580448 66728
rect 580500 66716 580506 66768
rect 66162 66648 66168 66700
rect 66220 66688 66226 66700
rect 187694 66688 187700 66700
rect 66220 66660 187700 66688
rect 66220 66648 66226 66660
rect 187694 66648 187700 66660
rect 187752 66648 187758 66700
rect 329098 66648 329104 66700
rect 329156 66688 329162 66700
rect 573358 66688 573364 66700
rect 329156 66660 573364 66688
rect 329156 66648 329162 66660
rect 573358 66648 573364 66660
rect 573416 66648 573422 66700
rect 68186 66580 68192 66632
rect 68244 66620 68250 66632
rect 168374 66620 168380 66632
rect 68244 66592 168380 66620
rect 68244 66580 68250 66592
rect 168374 66580 168380 66592
rect 168432 66580 168438 66632
rect 3418 66512 3424 66564
rect 3476 66552 3482 66564
rect 376570 66552 376576 66564
rect 3476 66524 376576 66552
rect 3476 66512 3482 66524
rect 376570 66512 376576 66524
rect 376628 66512 376634 66564
rect 3602 66172 3608 66224
rect 3660 66212 3666 66224
rect 90726 66212 90732 66224
rect 3660 66184 90732 66212
rect 3660 66172 3666 66184
rect 90726 66172 90732 66184
rect 90784 66172 90790 66224
rect 91002 66172 91008 66224
rect 91060 66212 91066 66224
rect 381906 66212 381912 66224
rect 91060 66184 381912 66212
rect 91060 66172 91066 66184
rect 381906 66172 381912 66184
rect 381964 66172 381970 66224
rect 403066 66172 403072 66224
rect 403124 66212 403130 66224
rect 575014 66212 575020 66224
rect 403124 66184 575020 66212
rect 403124 66172 403130 66184
rect 575014 66172 575020 66184
rect 575072 66172 575078 66224
rect 32398 66104 32404 66156
rect 32456 66144 32462 66156
rect 360746 66144 360752 66156
rect 32456 66116 360752 66144
rect 32456 66104 32462 66116
rect 360746 66104 360752 66116
rect 360804 66104 360810 66156
rect 371878 66104 371884 66156
rect 371936 66144 371942 66156
rect 535178 66144 535184 66156
rect 371936 66116 535184 66144
rect 371936 66104 371942 66116
rect 535178 66104 535184 66116
rect 535236 66104 535242 66156
rect 53742 66036 53748 66088
rect 53800 66076 53806 66088
rect 75178 66076 75184 66088
rect 53800 66048 75184 66076
rect 53800 66036 53806 66048
rect 75178 66036 75184 66048
rect 75236 66036 75242 66088
rect 80514 66036 80520 66088
rect 80572 66076 80578 66088
rect 81342 66076 81348 66088
rect 80572 66048 81348 66076
rect 80572 66036 80578 66048
rect 81342 66036 81348 66048
rect 81400 66036 81406 66088
rect 81529 66079 81587 66085
rect 81529 66045 81541 66079
rect 81575 66076 81587 66079
rect 440050 66076 440056 66088
rect 81575 66048 440056 66076
rect 81575 66045 81587 66048
rect 81529 66039 81587 66045
rect 440050 66036 440056 66048
rect 440108 66036 440114 66088
rect 450722 66036 450728 66088
rect 450780 66076 450786 66088
rect 574738 66076 574744 66088
rect 450780 66048 574744 66076
rect 450780 66036 450786 66048
rect 574738 66036 574744 66048
rect 574796 66036 574802 66088
rect 50430 65968 50436 66020
rect 50488 66008 50494 66020
rect 107010 66008 107016 66020
rect 50488 65980 107016 66008
rect 50488 65968 50494 65980
rect 107010 65968 107016 65980
rect 107068 65968 107074 66020
rect 130378 65968 130384 66020
rect 130436 66008 130442 66020
rect 508866 66008 508872 66020
rect 130436 65980 508872 66008
rect 130436 65968 130442 65980
rect 508866 65968 508872 65980
rect 508924 65968 508930 66020
rect 19242 65900 19248 65952
rect 19300 65940 19306 65952
rect 397730 65940 397736 65952
rect 19300 65912 397736 65940
rect 19300 65900 19306 65912
rect 397730 65900 397736 65912
rect 397788 65900 397794 65952
rect 24762 65832 24768 65884
rect 24820 65872 24826 65884
rect 159266 65872 159272 65884
rect 24820 65844 159272 65872
rect 24820 65832 24826 65844
rect 159266 65832 159272 65844
rect 159324 65832 159330 65884
rect 159358 65832 159364 65884
rect 159416 65872 159422 65884
rect 165154 65872 165160 65884
rect 159416 65844 165160 65872
rect 159416 65832 159422 65844
rect 165154 65832 165160 65844
rect 165212 65832 165218 65884
rect 184198 65832 184204 65884
rect 184256 65872 184262 65884
rect 571610 65872 571616 65884
rect 184256 65844 571616 65872
rect 184256 65832 184262 65844
rect 571610 65832 571616 65844
rect 571668 65832 571674 65884
rect 51718 65764 51724 65816
rect 51776 65804 51782 65816
rect 461210 65804 461216 65816
rect 51776 65776 461216 65804
rect 51776 65764 51782 65776
rect 461210 65764 461216 65776
rect 461268 65764 461274 65816
rect 60642 65696 60648 65748
rect 60700 65736 60706 65748
rect 85850 65736 85856 65748
rect 60700 65708 85856 65736
rect 60700 65696 60706 65708
rect 85850 65696 85856 65708
rect 85908 65696 85914 65748
rect 95142 65696 95148 65748
rect 95200 65736 95206 65748
rect 540514 65736 540520 65748
rect 95200 65708 540520 65736
rect 95200 65696 95206 65708
rect 540514 65696 540520 65708
rect 540572 65696 540578 65748
rect 53098 65628 53104 65680
rect 53156 65668 53162 65680
rect 498194 65668 498200 65680
rect 53156 65640 498200 65668
rect 53156 65628 53162 65640
rect 498194 65628 498200 65640
rect 498252 65628 498258 65680
rect 29638 65560 29644 65612
rect 29696 65600 29702 65612
rect 487706 65600 487712 65612
rect 29696 65572 487712 65600
rect 29696 65560 29702 65572
rect 487706 65560 487712 65572
rect 487764 65560 487770 65612
rect 47578 65492 47584 65544
rect 47636 65532 47642 65544
rect 567010 65532 567016 65544
rect 47636 65504 567016 65532
rect 47636 65492 47642 65504
rect 567010 65492 567016 65504
rect 567068 65492 567074 65544
rect 40678 65424 40684 65476
rect 40736 65464 40742 65476
rect 323762 65464 323768 65476
rect 40736 65436 323768 65464
rect 40736 65424 40742 65436
rect 323762 65424 323768 65436
rect 323820 65424 323826 65476
rect 345658 65424 345664 65476
rect 345716 65464 345722 65476
rect 355410 65464 355416 65476
rect 345716 65436 355416 65464
rect 345716 65424 345722 65436
rect 355410 65424 355416 65436
rect 355468 65424 355474 65476
rect 79318 65356 79324 65408
rect 79376 65396 79382 65408
rect 344922 65396 344928 65408
rect 79376 65368 344928 65396
rect 79376 65356 79382 65368
rect 344922 65356 344928 65368
rect 344980 65356 344986 65408
rect 28902 65288 28908 65340
rect 28960 65328 28966 65340
rect 133322 65328 133328 65340
rect 28960 65300 133328 65328
rect 28960 65288 28966 65300
rect 133322 65288 133328 65300
rect 133380 65288 133386 65340
rect 143994 65288 144000 65340
rect 144052 65328 144058 65340
rect 144822 65328 144828 65340
rect 144052 65300 144828 65328
rect 144052 65288 144058 65300
rect 144822 65288 144828 65300
rect 144880 65288 144886 65340
rect 160738 65288 160744 65340
rect 160796 65328 160802 65340
rect 424226 65328 424232 65340
rect 160796 65300 424232 65328
rect 160796 65288 160802 65300
rect 424226 65288 424232 65300
rect 424284 65288 424290 65340
rect 17862 65220 17868 65272
rect 17920 65260 17926 65272
rect 217962 65260 217968 65272
rect 17920 65232 217968 65260
rect 17920 65220 17926 65232
rect 217962 65220 217968 65232
rect 218020 65220 218026 65272
rect 235810 65220 235816 65272
rect 235868 65260 235874 65272
rect 276106 65260 276112 65272
rect 235868 65232 276112 65260
rect 235868 65220 235874 65232
rect 276106 65220 276112 65232
rect 276164 65220 276170 65272
rect 276658 65220 276664 65272
rect 276716 65260 276722 65272
rect 524690 65260 524696 65272
rect 276716 65232 524696 65260
rect 276716 65220 276722 65232
rect 524690 65220 524696 65232
rect 524748 65220 524754 65272
rect 33778 65152 33784 65204
rect 33836 65192 33842 65204
rect 228634 65192 228640 65204
rect 33836 65164 228640 65192
rect 33836 65152 33842 65164
rect 228634 65152 228640 65164
rect 228692 65152 228698 65204
rect 280798 65152 280804 65204
rect 280856 65192 280862 65204
rect 392578 65192 392584 65204
rect 280856 65164 392584 65192
rect 280856 65152 280862 65164
rect 392578 65152 392584 65164
rect 392636 65152 392642 65204
rect 35158 65084 35164 65136
rect 35216 65124 35222 65136
rect 191466 65124 191472 65136
rect 35216 65096 191472 65124
rect 35216 65084 35222 65096
rect 191466 65084 191472 65096
rect 191524 65084 191530 65136
rect 224862 65084 224868 65136
rect 224920 65124 224926 65136
rect 408402 65124 408408 65136
rect 224920 65096 408408 65124
rect 224920 65084 224926 65096
rect 408402 65084 408408 65096
rect 408460 65084 408466 65136
rect 70026 65016 70032 65068
rect 70084 65056 70090 65068
rect 81434 65056 81440 65068
rect 70084 65028 81440 65056
rect 70084 65016 70090 65028
rect 81434 65016 81440 65028
rect 81492 65016 81498 65068
rect 100662 65016 100668 65068
rect 100720 65056 100726 65068
rect 154482 65056 154488 65068
rect 100720 65028 154488 65056
rect 100720 65016 100726 65028
rect 154482 65016 154488 65028
rect 154540 65016 154546 65068
rect 181438 65016 181444 65068
rect 181496 65056 181502 65068
rect 281442 65056 281448 65068
rect 181496 65028 281448 65056
rect 181496 65016 181502 65028
rect 281442 65016 281448 65028
rect 281500 65016 281506 65068
rect 286318 65016 286324 65068
rect 286376 65056 286382 65068
rect 292114 65056 292120 65068
rect 286376 65028 292120 65056
rect 286376 65016 286382 65028
rect 292114 65016 292120 65028
rect 292172 65016 292178 65068
rect 297358 65016 297364 65068
rect 297416 65056 297422 65068
rect 371418 65056 371424 65068
rect 297416 65028 371424 65056
rect 297416 65016 297422 65028
rect 371418 65016 371424 65028
rect 371476 65016 371482 65068
rect 79962 64948 79968 65000
rect 80020 64988 80026 65000
rect 81529 64991 81587 64997
rect 81529 64988 81541 64991
rect 80020 64960 81541 64988
rect 80020 64948 80026 64960
rect 81529 64957 81541 64960
rect 81575 64957 81587 64991
rect 81529 64951 81587 64957
rect 104802 64948 104808 65000
rect 104860 64988 104866 65000
rect 112162 64988 112168 65000
rect 104860 64960 112168 64988
rect 104860 64948 104866 64960
rect 112162 64948 112168 64960
rect 112220 64948 112226 65000
rect 113082 64948 113088 65000
rect 113140 64988 113146 65000
rect 196802 64988 196808 65000
rect 113140 64960 196808 64988
rect 113140 64948 113146 64960
rect 196802 64948 196808 64960
rect 196860 64948 196866 65000
rect 291838 64948 291844 65000
rect 291896 64988 291902 65000
rect 318426 64988 318432 65000
rect 291896 64960 318432 64988
rect 291896 64948 291902 64960
rect 318426 64948 318432 64960
rect 318484 64948 318490 65000
rect 68462 64336 68468 64388
rect 68520 64376 68526 64388
rect 128354 64376 128360 64388
rect 68520 64348 128360 64376
rect 68520 64336 68526 64348
rect 128354 64336 128360 64348
rect 128412 64336 128418 64388
rect 138014 64336 138020 64388
rect 138072 64376 138078 64388
rect 162854 64376 162860 64388
rect 138072 64348 162860 64376
rect 138072 64336 138078 64348
rect 162854 64336 162860 64348
rect 162912 64336 162918 64388
rect 197262 64336 197268 64388
rect 197320 64376 197326 64388
rect 238754 64376 238760 64388
rect 197320 64348 238760 64376
rect 197320 64336 197326 64348
rect 238754 64336 238760 64348
rect 238812 64336 238818 64388
rect 117314 64268 117320 64320
rect 117372 64308 117378 64320
rect 230474 64308 230480 64320
rect 117372 64280 230480 64308
rect 117372 64268 117378 64280
rect 230474 64268 230480 64280
rect 230532 64268 230538 64320
rect 71038 64200 71044 64252
rect 71096 64240 71102 64252
rect 296714 64240 296720 64252
rect 71096 64212 296720 64240
rect 71096 64200 71102 64212
rect 296714 64200 296720 64212
rect 296772 64200 296778 64252
rect 122742 64132 122748 64184
rect 122800 64172 122806 64184
rect 569494 64172 569500 64184
rect 122800 64144 569500 64172
rect 122800 64132 122806 64144
rect 569494 64132 569500 64144
rect 569552 64132 569558 64184
rect 65518 62772 65524 62824
rect 65576 62812 65582 62824
rect 158714 62812 158720 62824
rect 65576 62784 158720 62812
rect 65576 62772 65582 62784
rect 158714 62772 158720 62784
rect 158772 62772 158778 62824
rect 194502 62772 194508 62824
rect 194560 62812 194566 62824
rect 572714 62812 572720 62824
rect 194560 62784 572720 62812
rect 194560 62772 194566 62784
rect 572714 62772 572720 62784
rect 572772 62772 572778 62824
rect 573450 60664 573456 60716
rect 573508 60704 573514 60716
rect 580166 60704 580172 60716
rect 573508 60676 580172 60704
rect 573508 60664 573514 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 11790 59344 11796 59356
rect 3108 59316 11796 59344
rect 3108 59304 3114 59316
rect 11790 59304 11796 59316
rect 11848 59304 11854 59356
rect 68278 57196 68284 57248
rect 68336 57236 68342 57248
rect 175274 57236 175280 57248
rect 68336 57208 175280 57236
rect 68336 57196 68342 57208
rect 175274 57196 175280 57208
rect 175332 57196 175338 57248
rect 67542 55836 67548 55888
rect 67600 55876 67606 55888
rect 580350 55876 580356 55888
rect 67600 55848 580356 55876
rect 67600 55836 67606 55848
rect 580350 55836 580356 55848
rect 580408 55836 580414 55888
rect 202690 46180 202696 46232
rect 202748 46220 202754 46232
rect 567746 46220 567752 46232
rect 202748 46192 567752 46220
rect 202748 46180 202754 46192
rect 567746 46180 567752 46192
rect 567804 46180 567810 46232
rect 59262 44140 59268 44192
rect 59320 44180 59326 44192
rect 64138 44180 64144 44192
rect 59320 44152 64144 44180
rect 59320 44140 59326 44152
rect 64138 44140 64144 44152
rect 64196 44140 64202 44192
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 149054 20652 149060 20664
rect 3476 20624 149060 20652
rect 3476 20612 3482 20624
rect 149054 20612 149060 20624
rect 149112 20612 149118 20664
rect 202782 20612 202788 20664
rect 202840 20652 202846 20664
rect 580166 20652 580172 20664
rect 202840 20624 580172 20652
rect 202840 20612 202846 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 144730 18572 144736 18624
rect 144788 18612 144794 18624
rect 249794 18612 249800 18624
rect 144788 18584 249800 18612
rect 144788 18572 144794 18584
rect 249794 18572 249800 18584
rect 249852 18572 249858 18624
rect 168374 11704 168380 11756
rect 168432 11744 168438 11756
rect 169570 11744 169576 11756
rect 168432 11716 169576 11744
rect 168432 11704 168438 11716
rect 169570 11704 169576 11716
rect 169628 11704 169634 11756
rect 71682 7760 71688 7812
rect 71740 7800 71746 7812
rect 311894 7800 311900 7812
rect 71740 7772 311900 7800
rect 71740 7760 71746 7772
rect 311894 7760 311900 7772
rect 311952 7760 311958 7812
rect 216858 7692 216864 7744
rect 216916 7732 216922 7744
rect 470594 7732 470600 7744
rect 216916 7704 470600 7732
rect 216916 7692 216922 7704
rect 470594 7692 470600 7704
rect 470652 7692 470658 7744
rect 131758 7624 131764 7676
rect 131816 7664 131822 7676
rect 429194 7664 429200 7676
rect 131816 7636 429200 7664
rect 131816 7624 131822 7636
rect 429194 7624 429200 7636
rect 429252 7624 429258 7676
rect 77386 7556 77392 7608
rect 77444 7596 77450 7608
rect 568574 7596 568580 7608
rect 77444 7568 568580 7596
rect 77444 7556 77450 7568
rect 568574 7556 568580 7568
rect 568632 7556 568638 7608
rect 134150 6808 134156 6860
rect 134208 6848 134214 6860
rect 244274 6848 244280 6860
rect 134208 6820 244280 6848
rect 134208 6808 134214 6820
rect 244274 6808 244280 6820
rect 244332 6808 244338 6860
rect 176654 6740 176660 6792
rect 176712 6780 176718 6792
rect 333974 6780 333980 6792
rect 176712 6752 333980 6780
rect 176712 6740 176718 6752
rect 333974 6740 333980 6752
rect 334032 6740 334038 6792
rect 192018 6672 192024 6724
rect 192076 6712 192082 6724
rect 349154 6712 349160 6724
rect 192076 6684 349160 6712
rect 192076 6672 192082 6684
rect 349154 6672 349160 6684
rect 349212 6672 349218 6724
rect 181530 6604 181536 6656
rect 181588 6644 181594 6656
rect 339494 6644 339500 6656
rect 181588 6616 339500 6644
rect 181588 6604 181594 6616
rect 339494 6604 339500 6616
rect 339552 6604 339558 6656
rect 142430 6536 142436 6588
rect 142488 6576 142494 6588
rect 160738 6576 160744 6588
rect 142488 6548 160744 6576
rect 142488 6536 142494 6548
rect 160738 6536 160744 6548
rect 160796 6536 160802 6588
rect 174262 6536 174268 6588
rect 174320 6576 174326 6588
rect 345658 6576 345664 6588
rect 174320 6548 345664 6576
rect 174320 6536 174326 6548
rect 345658 6536 345664 6548
rect 345716 6536 345722 6588
rect 138842 6468 138848 6520
rect 138900 6508 138906 6520
rect 159358 6508 159364 6520
rect 138900 6480 159364 6508
rect 138900 6468 138906 6480
rect 159358 6468 159364 6480
rect 159416 6468 159422 6520
rect 186130 6468 186136 6520
rect 186188 6508 186194 6520
rect 371878 6508 371884 6520
rect 186188 6480 371884 6508
rect 186188 6468 186194 6480
rect 371878 6468 371884 6480
rect 371936 6468 371942 6520
rect 148318 6400 148324 6452
rect 148376 6440 148382 6452
rect 434714 6440 434720 6452
rect 148376 6412 434720 6440
rect 148376 6400 148382 6412
rect 434714 6400 434720 6412
rect 434772 6400 434778 6452
rect 155402 6332 155408 6384
rect 155460 6372 155466 6384
rect 466454 6372 466460 6384
rect 155460 6344 466460 6372
rect 155460 6332 155466 6344
rect 466454 6332 466460 6344
rect 466512 6332 466518 6384
rect 144822 6264 144828 6316
rect 144880 6304 144886 6316
rect 173158 6304 173164 6316
rect 144880 6276 173164 6304
rect 144880 6264 144886 6276
rect 173158 6264 173164 6276
rect 173216 6264 173222 6316
rect 219250 6264 219256 6316
rect 219308 6304 219314 6316
rect 572898 6304 572904 6316
rect 219308 6276 572904 6304
rect 219308 6264 219314 6276
rect 572898 6264 572904 6276
rect 572956 6264 572962 6316
rect 147122 6196 147128 6248
rect 147180 6236 147186 6248
rect 518894 6236 518900 6248
rect 147180 6208 518900 6236
rect 147180 6196 147186 6208
rect 518894 6196 518900 6208
rect 518952 6196 518958 6248
rect 101030 6128 101036 6180
rect 101088 6168 101094 6180
rect 181438 6168 181444 6180
rect 101088 6140 181444 6168
rect 101088 6128 101094 6140
rect 181438 6128 181444 6140
rect 181496 6128 181502 6180
rect 187326 6128 187332 6180
rect 187384 6168 187390 6180
rect 572806 6168 572812 6180
rect 187384 6140 572812 6168
rect 187384 6128 187390 6140
rect 572806 6128 572812 6140
rect 572864 6128 572870 6180
rect 81342 5312 81348 5364
rect 81400 5352 81406 5364
rect 128170 5352 128176 5364
rect 81400 5324 128176 5352
rect 81400 5312 81406 5324
rect 128170 5312 128176 5324
rect 128228 5312 128234 5364
rect 69106 5244 69112 5296
rect 69164 5284 69170 5296
rect 96246 5284 96252 5296
rect 69164 5256 96252 5284
rect 69164 5244 69170 5256
rect 96246 5244 96252 5256
rect 96304 5244 96310 5296
rect 96522 5244 96528 5296
rect 96580 5284 96586 5296
rect 193214 5284 193220 5296
rect 96580 5256 193220 5284
rect 96580 5244 96586 5256
rect 193214 5244 193220 5256
rect 193272 5244 193278 5296
rect 232222 5244 232228 5296
rect 232280 5284 232286 5296
rect 412634 5284 412640 5296
rect 232280 5256 412640 5284
rect 232280 5244 232286 5256
rect 412634 5244 412640 5256
rect 412692 5244 412698 5296
rect 86862 5176 86868 5228
rect 86920 5216 86926 5228
rect 285674 5216 285680 5228
rect 86920 5188 285680 5216
rect 86920 5176 86926 5188
rect 285674 5176 285680 5188
rect 285732 5176 285738 5228
rect 31294 5108 31300 5160
rect 31352 5148 31358 5160
rect 270494 5148 270500 5160
rect 31352 5120 270500 5148
rect 31352 5108 31358 5120
rect 270494 5108 270500 5120
rect 270552 5108 270558 5160
rect 68094 5040 68100 5092
rect 68152 5080 68158 5092
rect 214466 5080 214472 5092
rect 68152 5052 214472 5080
rect 68152 5040 68158 5052
rect 214466 5040 214472 5052
rect 214524 5040 214530 5092
rect 235902 5040 235908 5092
rect 235960 5080 235966 5092
rect 481634 5080 481640 5092
rect 235960 5052 481640 5080
rect 235960 5040 235966 5052
rect 481634 5040 481640 5052
rect 481692 5040 481698 5092
rect 68646 4972 68652 5024
rect 68704 5012 68710 5024
rect 171962 5012 171968 5024
rect 68704 4984 171968 5012
rect 68704 4972 68710 4984
rect 171962 4972 171968 4984
rect 172020 4972 172026 5024
rect 177850 4972 177856 5024
rect 177908 5012 177914 5024
rect 207014 5012 207020 5024
rect 177908 4984 207020 5012
rect 177908 4972 177914 4984
rect 207014 4972 207020 4984
rect 207072 4972 207078 5024
rect 207382 4972 207388 5024
rect 207440 5012 207446 5024
rect 455414 5012 455420 5024
rect 207440 4984 455420 5012
rect 207440 4972 207446 4984
rect 455414 4972 455420 4984
rect 455472 4972 455478 5024
rect 65610 4904 65616 4956
rect 65668 4944 65674 4956
rect 137646 4944 137652 4956
rect 65668 4916 137652 4944
rect 65668 4904 65674 4916
rect 137646 4904 137652 4916
rect 137704 4904 137710 4956
rect 143534 4904 143540 4956
rect 143592 4944 143598 4956
rect 550634 4944 550640 4956
rect 143592 4916 550640 4944
rect 143592 4904 143598 4916
rect 550634 4904 550640 4916
rect 550692 4904 550698 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 130378 4876 130384 4888
rect 624 4848 130384 4876
rect 624 4836 630 4848
rect 130378 4836 130384 4848
rect 130436 4836 130442 4888
rect 136450 4836 136456 4888
rect 136508 4876 136514 4888
rect 572990 4876 572996 4888
rect 136508 4848 572996 4876
rect 136508 4836 136514 4848
rect 572990 4836 572996 4848
rect 573048 4836 573054 4888
rect 66714 4768 66720 4820
rect 66772 4808 66778 4820
rect 568942 4808 568948 4820
rect 66772 4780 568948 4808
rect 66772 4768 66778 4780
rect 568942 4768 568948 4780
rect 569000 4768 569006 4820
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 7650 4128 7656 4140
rect 6512 4100 7656 4128
rect 6512 4088 6518 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 69474 4020 69480 4072
rect 69532 4060 69538 4072
rect 98638 4060 98644 4072
rect 69532 4032 98644 4060
rect 69532 4020 69538 4032
rect 98638 4020 98644 4032
rect 98696 4020 98702 4072
rect 114002 4020 114008 4072
rect 114060 4060 114066 4072
rect 286318 4060 286324 4072
rect 114060 4032 286324 4060
rect 114060 4020 114066 4032
rect 286318 4020 286324 4032
rect 286376 4020 286382 4072
rect 64322 3952 64328 4004
rect 64380 3992 64386 4004
rect 276658 3992 276664 4004
rect 64380 3964 276664 3992
rect 64380 3952 64386 3964
rect 276658 3952 276664 3964
rect 276716 3952 276722 4004
rect 32490 3884 32496 3936
rect 32548 3924 32554 3936
rect 291838 3924 291844 3936
rect 32548 3896 291844 3924
rect 32548 3884 32554 3896
rect 291838 3884 291844 3896
rect 291896 3884 291902 3936
rect 14734 3816 14740 3868
rect 14792 3856 14798 3868
rect 280798 3856 280804 3868
rect 14792 3828 280804 3856
rect 14792 3816 14798 3828
rect 280798 3816 280804 3828
rect 280856 3816 280862 3868
rect 20622 3748 20628 3800
rect 20680 3788 20686 3800
rect 297358 3788 297364 3800
rect 20680 3760 297364 3788
rect 20680 3748 20686 3760
rect 297358 3748 297364 3760
rect 297416 3748 297422 3800
rect 44266 3680 44272 3732
rect 44324 3720 44330 3732
rect 47578 3720 47584 3732
rect 44324 3692 47584 3720
rect 44324 3680 44330 3692
rect 47578 3680 47584 3692
rect 47636 3680 47642 3732
rect 69750 3680 69756 3732
rect 69808 3720 69814 3732
rect 121086 3720 121092 3732
rect 69808 3692 121092 3720
rect 69808 3680 69814 3692
rect 121086 3680 121092 3692
rect 121144 3680 121150 3732
rect 215662 3680 215668 3732
rect 215720 3720 215726 3732
rect 568850 3720 568856 3732
rect 215720 3692 568856 3720
rect 215720 3680 215726 3692
rect 568850 3680 568856 3692
rect 568908 3680 568914 3732
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 22738 3652 22744 3664
rect 15988 3624 22744 3652
rect 15988 3612 15994 3624
rect 22738 3612 22744 3624
rect 22796 3612 22802 3664
rect 23014 3612 23020 3664
rect 23072 3652 23078 3664
rect 29638 3652 29644 3664
rect 23072 3624 29644 3652
rect 23072 3612 23078 3624
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 53098 3652 53104 3664
rect 45526 3624 53104 3652
rect 45526 3596 45554 3624
rect 53098 3612 53104 3624
rect 53156 3612 53162 3664
rect 69842 3612 69848 3664
rect 69900 3652 69906 3664
rect 123478 3652 123484 3664
rect 69900 3624 123484 3652
rect 69900 3612 69906 3624
rect 123478 3612 123484 3624
rect 123536 3612 123542 3664
rect 124674 3612 124680 3664
rect 124732 3652 124738 3664
rect 184198 3652 184204 3664
rect 124732 3624 184204 3652
rect 124732 3612 124738 3624
rect 184198 3612 184204 3624
rect 184256 3612 184262 3664
rect 213362 3612 213368 3664
rect 213420 3652 213426 3664
rect 569770 3652 569776 3664
rect 213420 3624 569776 3652
rect 213420 3612 213426 3624
rect 569770 3612 569776 3624
rect 569828 3612 569834 3664
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 11698 3584 11704 3596
rect 4120 3556 11704 3584
rect 4120 3544 4126 3556
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12308 3556 16574 3584
rect 12308 3544 12314 3556
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12342 3516 12348 3528
rect 11204 3488 12348 3516
rect 11204 3476 11210 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 16546 3516 16574 3556
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17862 3584 17868 3596
rect 17092 3556 17868 3584
rect 17092 3544 17098 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 19242 3584 19248 3596
rect 18288 3556 19248 3584
rect 18288 3544 18294 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 26142 3584 26148 3596
rect 25372 3556 26148 3584
rect 25372 3544 25378 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 26878 3584 26884 3596
rect 26436 3556 26884 3584
rect 26436 3516 26464 3556
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 35158 3584 35164 3596
rect 33652 3556 35164 3584
rect 33652 3544 33658 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 45462 3544 45468 3596
rect 45520 3556 45554 3596
rect 45520 3544 45526 3556
rect 48958 3544 48964 3596
rect 49016 3584 49022 3596
rect 58618 3584 58624 3596
rect 49016 3556 58624 3584
rect 49016 3544 49022 3556
rect 58618 3544 58624 3556
rect 58676 3544 58682 3596
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 61930 3584 61936 3596
rect 60884 3556 61936 3584
rect 60884 3544 60890 3556
rect 61930 3544 61936 3556
rect 61988 3544 61994 3596
rect 72418 3544 72424 3596
rect 72476 3584 72482 3596
rect 73985 3587 74043 3593
rect 72476 3556 73936 3584
rect 72476 3544 72482 3556
rect 16546 3488 26464 3516
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28902 3516 28908 3528
rect 27764 3488 28908 3516
rect 27764 3476 27770 3488
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 30098 3476 30104 3528
rect 30156 3516 30162 3528
rect 32398 3516 32404 3528
rect 30156 3488 32404 3516
rect 30156 3476 30162 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 39390 3516 39396 3528
rect 38436 3488 39396 3516
rect 38436 3476 38442 3488
rect 39390 3476 39396 3488
rect 39448 3476 39454 3528
rect 39574 3476 39580 3528
rect 39632 3516 39638 3528
rect 40678 3516 40684 3528
rect 39632 3488 40684 3516
rect 39632 3476 39638 3488
rect 40678 3476 40684 3488
rect 40736 3476 40742 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52362 3516 52368 3528
rect 51408 3488 52368 3516
rect 51408 3476 51414 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 57146 3516 57152 3528
rect 56100 3488 57152 3516
rect 56100 3476 56106 3488
rect 57146 3476 57152 3488
rect 57204 3476 57210 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 70302 3476 70308 3528
rect 70360 3516 70366 3528
rect 71038 3516 71044 3528
rect 70360 3488 71044 3516
rect 70360 3476 70366 3488
rect 71038 3476 71044 3488
rect 71096 3476 71102 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 73154 3476 73160 3528
rect 73212 3516 73218 3528
rect 73798 3516 73804 3528
rect 73212 3488 73804 3516
rect 73212 3476 73218 3488
rect 73798 3476 73804 3488
rect 73856 3476 73862 3528
rect 73908 3516 73936 3556
rect 73985 3553 73997 3587
rect 74031 3584 74043 3587
rect 94961 3587 95019 3593
rect 94961 3584 94973 3587
rect 74031 3556 94973 3584
rect 74031 3553 74043 3556
rect 73985 3547 74043 3553
rect 94961 3553 94973 3556
rect 95007 3553 95019 3587
rect 94961 3547 95019 3553
rect 95050 3544 95056 3596
rect 95108 3584 95114 3596
rect 95108 3556 103514 3584
rect 95108 3544 95114 3556
rect 89162 3516 89168 3528
rect 73908 3488 89168 3516
rect 89162 3476 89168 3488
rect 89220 3476 89226 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95142 3516 95148 3528
rect 94004 3488 95148 3516
rect 94004 3476 94010 3488
rect 95142 3476 95148 3488
rect 95200 3476 95206 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 103486 3516 103514 3556
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 115842 3584 115848 3596
rect 115256 3556 115848 3584
rect 115256 3544 115262 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 116394 3544 116400 3596
rect 116452 3584 116458 3596
rect 567838 3584 567844 3596
rect 116452 3556 567844 3584
rect 116452 3544 116458 3556
rect 567838 3544 567844 3556
rect 567896 3544 567902 3596
rect 570782 3516 570788 3528
rect 103486 3488 570788 3516
rect 570782 3476 570788 3488
rect 570840 3476 570846 3528
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 39298 3448 39304 3460
rect 1728 3420 39304 3448
rect 1728 3408 1734 3420
rect 39298 3408 39304 3420
rect 39356 3408 39362 3460
rect 51718 3448 51724 3460
rect 40696 3420 51724 3448
rect 40696 3392 40724 3420
rect 51718 3408 51724 3420
rect 51776 3408 51782 3460
rect 59630 3408 59636 3460
rect 59688 3448 59694 3460
rect 60642 3448 60648 3460
rect 59688 3420 60648 3448
rect 59688 3408 59694 3420
rect 60642 3408 60648 3420
rect 60700 3408 60706 3460
rect 69566 3408 69572 3460
rect 69624 3448 69630 3460
rect 73985 3451 74043 3457
rect 73985 3448 73997 3451
rect 69624 3420 73997 3448
rect 69624 3408 69630 3420
rect 73985 3417 73997 3420
rect 74031 3417 74043 3451
rect 85666 3448 85672 3460
rect 73985 3411 74043 3417
rect 74506 3420 85672 3448
rect 40678 3340 40684 3392
rect 40736 3340 40742 3392
rect 65886 3340 65892 3392
rect 65944 3380 65950 3392
rect 74506 3380 74534 3420
rect 85666 3408 85672 3420
rect 85724 3408 85730 3460
rect 87966 3408 87972 3460
rect 88024 3448 88030 3460
rect 569218 3448 569224 3460
rect 88024 3420 569224 3448
rect 88024 3408 88030 3420
rect 569218 3408 569224 3420
rect 569276 3408 569282 3460
rect 65944 3352 74534 3380
rect 65944 3340 65950 3352
rect 76190 3340 76196 3392
rect 76248 3380 76254 3392
rect 77202 3380 77208 3392
rect 76248 3352 77208 3380
rect 76248 3340 76254 3352
rect 77202 3340 77208 3352
rect 77260 3340 77266 3392
rect 78582 3340 78588 3392
rect 78640 3380 78646 3392
rect 79318 3380 79324 3392
rect 78640 3352 79324 3380
rect 78640 3340 78646 3352
rect 79318 3340 79324 3352
rect 79376 3340 79382 3392
rect 80146 3340 80152 3392
rect 80204 3380 80210 3392
rect 80882 3380 80888 3392
rect 80204 3352 80888 3380
rect 80204 3340 80210 3352
rect 80882 3340 80888 3352
rect 80940 3340 80946 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 94961 3383 95019 3389
rect 94961 3349 94973 3383
rect 95007 3380 95019 3383
rect 102226 3380 102232 3392
rect 95007 3352 102232 3380
rect 95007 3349 95019 3352
rect 94961 3343 95019 3349
rect 102226 3340 102232 3352
rect 102284 3340 102290 3392
rect 122282 3340 122288 3392
rect 122340 3380 122346 3392
rect 122742 3380 122748 3392
rect 122340 3352 122748 3380
rect 122340 3340 122346 3352
rect 122742 3340 122748 3352
rect 122800 3340 122806 3392
rect 125870 3340 125876 3392
rect 125928 3380 125934 3392
rect 126882 3380 126888 3392
rect 125928 3352 126888 3380
rect 125928 3340 125934 3352
rect 126882 3340 126888 3352
rect 126940 3340 126946 3392
rect 126974 3340 126980 3392
rect 127032 3380 127038 3392
rect 128262 3380 128268 3392
rect 127032 3352 128268 3380
rect 127032 3340 127038 3352
rect 128262 3340 128268 3352
rect 128320 3340 128326 3392
rect 149514 3340 149520 3392
rect 149572 3380 149578 3392
rect 150342 3380 150348 3392
rect 149572 3352 150348 3380
rect 149572 3340 149578 3352
rect 150342 3340 150348 3352
rect 150400 3340 150406 3392
rect 151814 3340 151820 3392
rect 151872 3380 151878 3392
rect 153102 3380 153108 3392
rect 151872 3352 153108 3380
rect 151872 3340 151878 3352
rect 153102 3340 153108 3352
rect 153160 3340 153166 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186038 3380 186044 3392
rect 184992 3352 186044 3380
rect 184992 3340 184998 3352
rect 186038 3340 186044 3352
rect 186096 3340 186102 3392
rect 189718 3340 189724 3392
rect 189776 3380 189782 3392
rect 190362 3380 190368 3392
rect 189776 3352 190368 3380
rect 189776 3340 189782 3352
rect 190362 3340 190368 3352
rect 190420 3340 190426 3392
rect 196802 3340 196808 3392
rect 196860 3380 196866 3392
rect 197262 3380 197268 3392
rect 196860 3352 197268 3380
rect 196860 3340 196866 3352
rect 197262 3340 197268 3352
rect 197320 3340 197326 3392
rect 199102 3340 199108 3392
rect 199160 3380 199166 3392
rect 200022 3380 200028 3392
rect 199160 3352 200028 3380
rect 199160 3340 199166 3352
rect 200022 3340 200028 3352
rect 200080 3340 200086 3392
rect 206186 3340 206192 3392
rect 206244 3380 206250 3392
rect 206922 3380 206928 3392
rect 206244 3352 206928 3380
rect 206244 3340 206250 3352
rect 206922 3340 206928 3352
rect 206980 3340 206986 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219342 3380 219348 3392
rect 218112 3352 219348 3380
rect 218112 3340 218118 3352
rect 219342 3340 219348 3352
rect 219400 3340 219406 3392
rect 223942 3340 223948 3392
rect 224000 3380 224006 3392
rect 224862 3380 224868 3392
rect 224000 3352 224868 3380
rect 224000 3340 224006 3352
rect 224862 3340 224868 3352
rect 224920 3340 224926 3392
rect 225138 3340 225144 3392
rect 225196 3380 225202 3392
rect 226242 3380 226248 3392
rect 225196 3352 226248 3380
rect 225196 3340 225202 3352
rect 226242 3340 226248 3352
rect 226300 3340 226306 3392
rect 229830 3340 229836 3392
rect 229888 3380 229894 3392
rect 230382 3380 230388 3392
rect 229888 3352 230388 3380
rect 229888 3340 229894 3352
rect 230382 3340 230388 3352
rect 230440 3340 230446 3392
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 235810 3380 235816 3392
rect 234672 3352 235816 3380
rect 234672 3340 234678 3352
rect 235810 3340 235816 3352
rect 235868 3340 235874 3392
rect 28902 3204 28908 3256
rect 28960 3244 28966 3256
rect 33778 3244 33784 3256
rect 28960 3216 33784 3244
rect 28960 3204 28966 3216
rect 33778 3204 33784 3216
rect 33836 3204 33842 3256
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 4982 3176 4988 3188
rect 2924 3148 4988 3176
rect 2924 3136 2930 3148
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 10318 3176 10324 3188
rect 7708 3148 10324 3176
rect 7708 3136 7714 3148
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 21358 3040 21364 3052
rect 19484 3012 21364 3040
rect 19484 3000 19490 3012
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 47854 3000 47860 3052
rect 47912 3040 47918 3052
rect 50338 3040 50344 3052
rect 47912 3012 50344 3040
rect 47912 3000 47918 3012
rect 50338 3000 50344 3012
rect 50396 3000 50402 3052
rect 52546 3000 52552 3052
rect 52604 3040 52610 3052
rect 54478 3040 54484 3052
rect 52604 3012 54484 3040
rect 52604 3000 52610 3012
rect 54478 3000 54484 3012
rect 54536 3000 54542 3052
rect 69106 2932 69112 2984
rect 69164 2972 69170 2984
rect 71682 2972 71688 2984
rect 69164 2944 71688 2972
rect 69164 2932 69170 2944
rect 71682 2932 71688 2944
rect 71740 2932 71746 2984
rect 24210 2864 24216 2916
rect 24268 2904 24274 2916
rect 24762 2904 24768 2916
rect 24268 2876 24768 2904
rect 24268 2864 24274 2876
rect 24762 2864 24768 2876
rect 24820 2864 24826 2916
<< via1 >>
rect 283840 700816 283892 700868
rect 439596 700816 439648 700868
rect 318708 700748 318760 700800
rect 478512 700748 478564 700800
rect 170312 700680 170364 700732
rect 333980 700680 334032 700732
rect 348792 700680 348844 700732
rect 439504 700680 439556 700732
rect 154120 700612 154172 700664
rect 418160 700612 418212 700664
rect 300124 700544 300176 700596
rect 570328 700544 570380 700596
rect 277308 700476 277360 700528
rect 559656 700476 559708 700528
rect 69848 700408 69900 700460
rect 364984 700408 365036 700460
rect 413652 700408 413704 700460
rect 568856 700408 568908 700460
rect 89168 700340 89220 700392
rect 424324 700340 424376 700392
rect 543464 700340 543516 700392
rect 568580 700340 568632 700392
rect 40500 700272 40552 700324
rect 105544 700272 105596 700324
rect 218980 700272 219032 700324
rect 570052 700272 570104 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 494796 699660 494848 699712
rect 495348 699660 495400 699712
rect 3424 683136 3476 683188
rect 569960 683136 570012 683188
rect 576216 683136 576268 683188
rect 580172 683136 580224 683188
rect 2780 671032 2832 671084
rect 4804 671032 4856 671084
rect 573364 670692 573416 670744
rect 580172 670692 580224 670744
rect 3424 632068 3476 632120
rect 570420 632068 570472 632120
rect 68744 630640 68796 630692
rect 580172 630640 580224 630692
rect 256608 616836 256660 616888
rect 580172 616836 580224 616888
rect 2780 579912 2832 579964
rect 4896 579912 4948 579964
rect 574744 576852 574796 576904
rect 580172 576852 580224 576904
rect 105544 571276 105596 571328
rect 107200 571276 107252 571328
rect 276480 571276 276532 571328
rect 277308 571276 277360 571328
rect 64144 571004 64196 571056
rect 186504 571004 186556 571056
rect 10324 570936 10376 570988
rect 530216 570936 530268 570988
rect 58624 570800 58676 570852
rect 138848 570800 138900 570852
rect 57244 570732 57296 570784
rect 149520 570732 149572 570784
rect 255320 570732 255372 570784
rect 256608 570732 256660 570784
rect 439504 570732 439556 570784
rect 472072 570732 472124 570784
rect 495348 570732 495400 570784
rect 535552 570732 535604 570784
rect 54484 570664 54536 570716
rect 165344 570664 165396 570716
rect 439596 570664 439648 570716
rect 556712 570664 556764 570716
rect 12348 570596 12400 570648
rect 123024 570596 123076 570648
rect 424324 570596 424376 570648
rect 561864 570596 561916 570648
rect 65524 570528 65576 570580
rect 191840 570528 191892 570580
rect 68836 570460 68888 570512
rect 239312 570460 239364 570512
rect 22744 570392 22796 570444
rect 196992 570392 197044 570444
rect 178132 570324 178184 570376
rect 456248 570324 456300 570376
rect 39304 570256 39356 570308
rect 350448 570256 350500 570308
rect 408592 570256 408644 570308
rect 569316 570256 569368 570308
rect 50344 570188 50396 570240
rect 450912 570188 450964 570240
rect 69664 570120 69716 570172
rect 477408 570120 477460 570172
rect 66076 570052 66128 570104
rect 487896 570052 487948 570104
rect 26884 569984 26936 570036
rect 509056 569984 509108 570036
rect 68928 569916 68980 569968
rect 75368 569916 75420 569968
rect 234160 568216 234212 568268
rect 573456 568216 573508 568268
rect 11704 568148 11756 568200
rect 355784 568148 355836 568200
rect 10416 568080 10468 568132
rect 360936 568080 360988 568132
rect 398104 568080 398156 568132
rect 576308 568080 576360 568132
rect 5080 568012 5132 568064
rect 218336 568012 218388 568064
rect 223304 568012 223356 568064
rect 580264 568012 580316 568064
rect 7656 567944 7708 567996
rect 365996 567944 366048 567996
rect 371976 567944 372028 567996
rect 577504 567944 577556 567996
rect 208032 567876 208084 567928
rect 573548 567876 573600 567928
rect 46848 567808 46900 567860
rect 424140 567808 424192 567860
rect 3424 567740 3476 567792
rect 159732 567740 159784 567792
rect 202696 567740 202748 567792
rect 580356 567740 580408 567792
rect 44088 567672 44140 567724
rect 429476 567672 429528 567724
rect 11796 567604 11848 567656
rect 434812 567604 434864 567656
rect 445760 567604 445812 567656
rect 574928 567604 574980 567656
rect 62028 567536 62080 567588
rect 492956 567536 493008 567588
rect 118056 567468 118108 567520
rect 574836 567468 574888 567520
rect 112812 567400 112864 567452
rect 576124 567400 576176 567452
rect 39396 567332 39448 567384
rect 514116 567332 514168 567384
rect 66168 567264 66220 567316
rect 69940 567264 69992 567316
rect 91744 567264 91796 567316
rect 96712 567264 96764 567316
rect 571248 567264 571300 567316
rect 570604 567196 570656 567248
rect 3608 566448 3660 566500
rect 570236 566448 570288 566500
rect 3516 566312 3568 566364
rect 7564 566312 7616 566364
rect 568764 565972 568816 566024
rect 69020 565836 69072 565888
rect 568580 565904 568632 565956
rect 569408 565904 569460 565956
rect 571248 564340 571300 564392
rect 580172 564340 580224 564392
rect 68652 561688 68704 561740
rect 69020 561688 69072 561740
rect 4988 560260 5040 560312
rect 67640 560260 67692 560312
rect 64880 559852 64932 559904
rect 68652 559852 68704 559904
rect 57888 556180 57940 556232
rect 64788 556180 64840 556232
rect 571340 554752 571392 554804
rect 573732 554752 573784 554804
rect 55864 551760 55916 551812
rect 57888 551760 57940 551812
rect 568948 548088 569000 548140
rect 569408 548088 569460 548140
rect 47584 546388 47636 546440
rect 55864 546456 55916 546508
rect 568948 540379 569000 540388
rect 568948 540345 568957 540379
rect 568957 540345 568991 540379
rect 568991 540345 569000 540379
rect 568948 540336 569000 540345
rect 65984 536800 66036 536852
rect 67640 536800 67692 536852
rect 42064 532040 42116 532092
rect 47584 532040 47636 532092
rect 568948 525351 569000 525360
rect 568948 525317 568957 525351
rect 568957 525317 568991 525351
rect 568991 525317 569000 525351
rect 568948 525308 569000 525317
rect 39672 514768 39724 514820
rect 42064 514768 42116 514820
rect 571984 511912 572036 511964
rect 580172 511912 580224 511964
rect 37188 510552 37240 510604
rect 39672 510620 39724 510672
rect 568948 503047 569000 503056
rect 568948 503013 568957 503047
rect 568957 503013 568991 503047
rect 568991 503013 569000 503047
rect 568948 503004 569000 503013
rect 35164 502936 35216 502988
rect 37188 502936 37240 502988
rect 569040 499740 569092 499792
rect 569408 499740 569460 499792
rect 568948 498040 569000 498092
rect 568948 497904 569000 497956
rect 569408 497904 569460 497956
rect 568948 497768 569000 497820
rect 568948 495363 569000 495372
rect 568948 495329 568957 495363
rect 568957 495329 568991 495363
rect 568991 495329 569000 495363
rect 568948 495320 569000 495329
rect 33232 491240 33284 491292
rect 35164 491240 35216 491292
rect 32404 487160 32456 487212
rect 33232 487160 33284 487212
rect 568948 486455 569000 486464
rect 568948 486421 568957 486455
rect 568957 486421 568991 486455
rect 568991 486421 569000 486455
rect 568948 486412 569000 486421
rect 568948 485095 569000 485104
rect 568948 485061 568957 485095
rect 568957 485061 568991 485095
rect 568991 485061 569000 485095
rect 568948 485052 569000 485061
rect 30380 478864 30432 478916
rect 32404 478864 32456 478916
rect 571340 477640 571392 477692
rect 573640 477640 573692 477692
rect 2780 475872 2832 475924
rect 5080 475872 5132 475924
rect 25136 469820 25188 469872
rect 30012 469820 30064 469872
rect 24124 466420 24176 466472
rect 25136 466420 25188 466472
rect 570604 458124 570656 458176
rect 580172 458124 580224 458176
rect 68652 451120 68704 451172
rect 69756 451120 69808 451172
rect 568948 445748 569000 445800
rect 569408 445748 569460 445800
rect 568948 431536 569000 431588
rect 569408 431536 569460 431588
rect 65800 426436 65852 426488
rect 67916 426436 67968 426488
rect 22836 424736 22888 424788
rect 24124 424736 24176 424788
rect 2780 423512 2832 423564
rect 5080 423512 5132 423564
rect 575020 418140 575072 418192
rect 580172 418140 580224 418192
rect 21364 417324 21416 417376
rect 22836 417324 22888 417376
rect 13728 411272 13780 411324
rect 67640 411272 67692 411324
rect 3332 409844 3384 409896
rect 50436 409844 50488 409896
rect 18604 408756 18656 408808
rect 21364 408756 21416 408808
rect 15844 407192 15896 407244
rect 18604 407192 18656 407244
rect 573732 405628 573784 405680
rect 580172 405628 580224 405680
rect 65892 403248 65944 403300
rect 68008 403248 68060 403300
rect 12440 400188 12492 400240
rect 15844 400188 15896 400240
rect 5540 396720 5592 396772
rect 12440 396720 12492 396772
rect 3976 396040 4028 396092
rect 67640 396040 67692 396092
rect 569224 390532 569276 390584
rect 571708 390532 571760 390584
rect 3700 372580 3752 372632
rect 67640 372580 67692 372632
rect 3240 371220 3292 371272
rect 5172 371220 5224 371272
rect 569316 365644 569368 365696
rect 579988 365644 580040 365696
rect 55128 364352 55180 364404
rect 67640 364352 67692 364404
rect 65708 356056 65760 356108
rect 67824 356056 67876 356108
rect 3516 350480 3568 350532
rect 67640 350480 67692 350532
rect 572076 344972 572128 345024
rect 575020 344972 575072 345024
rect 52368 342864 52420 342916
rect 65524 342864 65576 342916
rect 572628 329536 572680 329588
rect 576216 329536 576268 329588
rect 24768 327020 24820 327072
rect 67640 327020 67692 327072
rect 568948 321580 569000 321632
rect 569316 321580 569368 321632
rect 3516 320084 3568 320136
rect 7656 320084 7708 320136
rect 68192 310428 68244 310480
rect 69848 310428 69900 310480
rect 571340 305600 571392 305652
rect 572996 305600 573048 305652
rect 27528 302880 27580 302932
rect 68284 302880 68336 302932
rect 65524 302200 65576 302252
rect 67824 302200 67876 302252
rect 576308 299412 576360 299464
rect 580172 299412 580224 299464
rect 65616 285676 65668 285728
rect 67824 285676 67876 285728
rect 3884 270512 3936 270564
rect 67640 270512 67692 270564
rect 569040 266364 569092 266416
rect 569316 266364 569368 266416
rect 569132 258476 569184 258528
rect 569316 258476 569368 258528
rect 575020 258068 575072 258120
rect 579620 258068 579672 258120
rect 68376 247664 68428 247716
rect 69848 247664 69900 247716
rect 574928 245556 574980 245608
rect 580172 245556 580224 245608
rect 63408 238756 63460 238808
rect 67640 238756 67692 238808
rect 10968 231820 11020 231872
rect 67640 231820 67692 231872
rect 568948 219716 569000 219768
rect 569408 219716 569460 219768
rect 574928 218016 574980 218068
rect 580172 218016 580224 218068
rect 26148 208360 26200 208412
rect 67640 208360 67692 208412
rect 68376 193128 68428 193180
rect 69572 193128 69624 193180
rect 3332 187688 3384 187740
rect 5172 187688 5224 187740
rect 577504 179324 577556 179376
rect 579896 179324 579948 179376
rect 9588 176672 9640 176724
rect 67640 176672 67692 176724
rect 5540 171096 5592 171148
rect 8300 171028 8352 171080
rect 8300 168376 8352 168428
rect 9772 168376 9824 168428
rect 574836 166948 574888 167000
rect 580172 166948 580224 167000
rect 9772 164228 9824 164280
rect 15200 164160 15252 164212
rect 65432 161508 65484 161560
rect 67640 161508 67692 161560
rect 15200 161372 15252 161424
rect 19248 161372 19300 161424
rect 19340 151784 19392 151836
rect 22836 151716 22888 151768
rect 2780 150084 2832 150136
rect 4988 150084 5040 150136
rect 68100 146208 68152 146260
rect 69480 146208 69532 146260
rect 570788 140768 570840 140820
rect 571800 140768 571852 140820
rect 3608 139340 3660 139392
rect 67640 139340 67692 139392
rect 573640 139340 573692 139392
rect 580172 139340 580224 139392
rect 22836 138660 22888 138712
rect 24124 138660 24176 138712
rect 24124 129752 24176 129804
rect 66812 129752 66864 129804
rect 67640 129752 67692 129804
rect 28264 129684 28316 129736
rect 573548 126896 573600 126948
rect 579620 126896 579672 126948
rect 28264 125536 28316 125588
rect 30288 125536 30340 125588
rect 30380 118124 30432 118176
rect 32404 118124 32456 118176
rect 32404 105476 32456 105528
rect 37280 105476 37332 105528
rect 37280 100852 37332 100904
rect 40040 100852 40092 100904
rect 576124 100648 576176 100700
rect 579712 100648 579764 100700
rect 22008 97996 22060 98048
rect 67640 97996 67692 98048
rect 3332 97928 3384 97980
rect 10416 97928 10468 97980
rect 40040 95140 40092 95192
rect 42616 95140 42668 95192
rect 42616 92284 42668 92336
rect 44180 92284 44232 92336
rect 44180 90312 44232 90364
rect 49608 90312 49660 90364
rect 49700 86912 49752 86964
rect 52276 86912 52328 86964
rect 37188 82832 37240 82884
rect 68376 82832 68428 82884
rect 52276 82424 52328 82476
rect 56508 82424 56560 82476
rect 569776 80044 569828 80096
rect 571524 80044 571576 80096
rect 56508 77256 56560 77308
rect 63500 77188 63552 77240
rect 63500 75148 63552 75200
rect 69388 75148 69440 75200
rect 569316 71136 569368 71188
rect 569868 71136 569920 71188
rect 50988 70048 51040 70100
rect 570604 70048 570656 70100
rect 42708 69980 42760 70032
rect 570328 69980 570380 70032
rect 37096 69912 37148 69964
rect 570512 69912 570564 69964
rect 35808 69844 35860 69896
rect 570972 69844 571024 69896
rect 21364 69776 21416 69828
rect 567844 69776 567896 69828
rect 571984 69776 572036 69828
rect 7656 69708 7708 69760
rect 572076 69708 572128 69760
rect 4988 69640 5040 69692
rect 571340 69640 571392 69692
rect 57888 69572 57940 69624
rect 571432 69572 571484 69624
rect 69020 69504 69072 69556
rect 580540 69504 580592 69556
rect 67640 69436 67692 69488
rect 580264 69436 580316 69488
rect 61936 69368 61988 69420
rect 572260 69368 572312 69420
rect 65340 69300 65392 69352
rect 569040 69300 569092 69352
rect 69388 69232 69440 69284
rect 569592 69232 569644 69284
rect 571892 69164 571944 69216
rect 68376 68960 68428 69012
rect 68744 69096 68796 69148
rect 68744 68960 68796 69012
rect 68928 68960 68980 69012
rect 569408 68960 569460 69012
rect 67732 68892 67784 68944
rect 570420 68892 570472 68944
rect 67916 68824 67968 68876
rect 569684 68824 569736 68876
rect 68928 68756 68980 68808
rect 69664 68756 69716 68808
rect 569960 68756 570012 68808
rect 66996 68688 67048 68740
rect 69296 68688 69348 68740
rect 70400 68688 70452 68740
rect 68560 68620 68612 68672
rect 132592 68688 132644 68740
rect 153108 68688 153160 68740
rect 572536 68688 572588 68740
rect 67824 68552 67876 68604
rect 72424 68552 72476 68604
rect 66812 68484 66864 68536
rect 140780 68620 140832 68672
rect 572444 68620 572496 68672
rect 128360 68552 128412 68604
rect 570236 68552 570288 68604
rect 84200 68484 84252 68536
rect 126888 68484 126940 68536
rect 570052 68484 570104 68536
rect 68836 68416 68888 68468
rect 80152 68416 80204 68468
rect 84108 68416 84160 68468
rect 568672 68416 568724 68468
rect 66076 68348 66128 68400
rect 73160 68348 73212 68400
rect 77208 68348 77260 68400
rect 569316 68348 569368 68400
rect 65708 68280 65760 68332
rect 73068 68280 73120 68332
rect 572168 68280 572220 68332
rect 66904 68212 66956 68264
rect 190552 68212 190604 68264
rect 197360 68255 197412 68264
rect 197360 68221 197369 68255
rect 197369 68221 197403 68255
rect 197403 68221 197412 68255
rect 197360 68212 197412 68221
rect 200028 68255 200080 68264
rect 200028 68221 200037 68255
rect 200037 68221 200071 68255
rect 200071 68221 200080 68255
rect 200028 68212 200080 68221
rect 206928 68212 206980 68264
rect 571800 68212 571852 68264
rect 67180 68144 67232 68196
rect 211160 68144 211212 68196
rect 219348 68144 219400 68196
rect 570696 68144 570748 68196
rect 67364 68076 67416 68128
rect 222200 68076 222252 68128
rect 226248 68076 226300 68128
rect 570144 68076 570196 68128
rect 68744 68008 68796 68060
rect 227812 68008 227864 68060
rect 230388 68008 230440 68060
rect 569132 68008 569184 68060
rect 69204 67940 69256 67992
rect 74632 67940 74684 67992
rect 220820 67940 220872 67992
rect 65800 67872 65852 67924
rect 209780 67872 209832 67924
rect 65432 67804 65484 67856
rect 167000 67804 167052 67856
rect 178040 67847 178092 67856
rect 178040 67813 178049 67847
rect 178049 67813 178083 67847
rect 178083 67813 178092 67847
rect 178040 67804 178092 67813
rect 182180 67847 182232 67856
rect 182180 67813 182189 67847
rect 182189 67813 182223 67847
rect 182223 67813 182232 67847
rect 182180 67804 182232 67813
rect 186044 67847 186096 67856
rect 186044 67813 186053 67847
rect 186053 67813 186087 67847
rect 186087 67813 186096 67847
rect 186044 67804 186096 67813
rect 190368 67847 190420 67856
rect 190368 67813 190377 67847
rect 190377 67813 190411 67847
rect 190411 67813 190420 67847
rect 190368 67804 190420 67813
rect 67272 67736 67324 67788
rect 161480 67736 161532 67788
rect 68008 67668 68060 67720
rect 157340 67668 157392 67720
rect 68376 67600 68428 67652
rect 150348 67600 150400 67652
rect 154304 67643 154356 67652
rect 154304 67609 154313 67643
rect 154313 67609 154347 67643
rect 154347 67609 154356 67643
rect 154304 67600 154356 67609
rect 4896 67532 4948 67584
rect 545856 67532 545908 67584
rect 4804 67464 4856 67516
rect 503536 67464 503588 67516
rect 4068 67396 4120 67448
rect 477040 67396 477092 67448
rect 7564 67328 7616 67380
rect 418896 67328 418948 67380
rect 3792 67260 3844 67312
rect 387248 67260 387300 67312
rect 5080 67192 5132 67244
rect 128176 67192 128228 67244
rect 366088 67192 366140 67244
rect 574928 67192 574980 67244
rect 119988 67124 120040 67176
rect 572352 67124 572404 67176
rect 115848 67056 115900 67108
rect 568764 67056 568816 67108
rect 65984 66988 66036 67040
rect 91100 66988 91152 67040
rect 111708 66988 111760 67040
rect 569868 66988 569920 67040
rect 67088 66920 67140 66972
rect 580264 66920 580316 66972
rect 3700 66852 3752 66904
rect 570880 66852 570932 66904
rect 3516 66784 3568 66836
rect 175648 66784 175700 66836
rect 254952 66784 255004 66836
rect 580356 66784 580408 66836
rect 67456 66716 67508 66768
rect 208400 66716 208452 66768
rect 260288 66716 260340 66768
rect 580448 66716 580500 66768
rect 66168 66648 66220 66700
rect 187700 66648 187752 66700
rect 329104 66648 329156 66700
rect 573364 66648 573416 66700
rect 68192 66580 68244 66632
rect 168380 66580 168432 66632
rect 3424 66512 3476 66564
rect 376576 66512 376628 66564
rect 3608 66172 3660 66224
rect 90732 66172 90784 66224
rect 91008 66172 91060 66224
rect 381912 66172 381964 66224
rect 403072 66172 403124 66224
rect 575020 66172 575072 66224
rect 32404 66104 32456 66156
rect 360752 66104 360804 66156
rect 371884 66104 371936 66156
rect 535184 66104 535236 66156
rect 53748 66036 53800 66088
rect 75184 66036 75236 66088
rect 80520 66036 80572 66088
rect 81348 66036 81400 66088
rect 440056 66036 440108 66088
rect 450728 66036 450780 66088
rect 574744 66036 574796 66088
rect 50436 65968 50488 66020
rect 107016 65968 107068 66020
rect 130384 65968 130436 66020
rect 508872 65968 508924 66020
rect 19248 65900 19300 65952
rect 397736 65900 397788 65952
rect 24768 65832 24820 65884
rect 159272 65832 159324 65884
rect 159364 65832 159416 65884
rect 165160 65832 165212 65884
rect 184204 65832 184256 65884
rect 571616 65832 571668 65884
rect 51724 65764 51776 65816
rect 461216 65764 461268 65816
rect 60648 65696 60700 65748
rect 85856 65696 85908 65748
rect 95148 65696 95200 65748
rect 540520 65696 540572 65748
rect 53104 65628 53156 65680
rect 498200 65628 498252 65680
rect 29644 65560 29696 65612
rect 487712 65560 487764 65612
rect 47584 65492 47636 65544
rect 567016 65492 567068 65544
rect 40684 65424 40736 65476
rect 323768 65424 323820 65476
rect 345664 65424 345716 65476
rect 355416 65424 355468 65476
rect 79324 65356 79376 65408
rect 344928 65356 344980 65408
rect 28908 65288 28960 65340
rect 133328 65288 133380 65340
rect 144000 65288 144052 65340
rect 144828 65288 144880 65340
rect 160744 65288 160796 65340
rect 424232 65288 424284 65340
rect 17868 65220 17920 65272
rect 217968 65220 218020 65272
rect 235816 65220 235868 65272
rect 276112 65220 276164 65272
rect 276664 65220 276716 65272
rect 524696 65220 524748 65272
rect 33784 65152 33836 65204
rect 228640 65152 228692 65204
rect 280804 65152 280856 65204
rect 392584 65152 392636 65204
rect 35164 65084 35216 65136
rect 191472 65084 191524 65136
rect 224868 65084 224920 65136
rect 408408 65084 408460 65136
rect 70032 65016 70084 65068
rect 81440 65016 81492 65068
rect 100668 65016 100720 65068
rect 154488 65016 154540 65068
rect 181444 65016 181496 65068
rect 281448 65016 281500 65068
rect 286324 65016 286376 65068
rect 292120 65016 292172 65068
rect 297364 65016 297416 65068
rect 371424 65016 371476 65068
rect 79968 64948 80020 65000
rect 104808 64948 104860 65000
rect 112168 64948 112220 65000
rect 113088 64948 113140 65000
rect 196808 64948 196860 65000
rect 291844 64948 291896 65000
rect 318432 64948 318484 65000
rect 68468 64336 68520 64388
rect 128360 64336 128412 64388
rect 138020 64336 138072 64388
rect 162860 64336 162912 64388
rect 197268 64336 197320 64388
rect 238760 64336 238812 64388
rect 117320 64268 117372 64320
rect 230480 64268 230532 64320
rect 71044 64200 71096 64252
rect 296720 64200 296772 64252
rect 122748 64132 122800 64184
rect 569500 64132 569552 64184
rect 65524 62772 65576 62824
rect 158720 62772 158772 62824
rect 194508 62772 194560 62824
rect 572720 62772 572772 62824
rect 573456 60664 573508 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 11796 59304 11848 59356
rect 68284 57196 68336 57248
rect 175280 57196 175332 57248
rect 67548 55836 67600 55888
rect 580356 55836 580408 55888
rect 202696 46180 202748 46232
rect 567752 46180 567804 46232
rect 59268 44140 59320 44192
rect 64144 44140 64196 44192
rect 3424 20612 3476 20664
rect 149060 20612 149112 20664
rect 202788 20612 202840 20664
rect 580172 20612 580224 20664
rect 144736 18572 144788 18624
rect 249800 18572 249852 18624
rect 168380 11704 168432 11756
rect 169576 11704 169628 11756
rect 71688 7760 71740 7812
rect 311900 7760 311952 7812
rect 216864 7692 216916 7744
rect 470600 7692 470652 7744
rect 131764 7624 131816 7676
rect 429200 7624 429252 7676
rect 77392 7556 77444 7608
rect 568580 7556 568632 7608
rect 134156 6808 134208 6860
rect 244280 6808 244332 6860
rect 176660 6740 176712 6792
rect 333980 6740 334032 6792
rect 192024 6672 192076 6724
rect 349160 6672 349212 6724
rect 181536 6604 181588 6656
rect 339500 6604 339552 6656
rect 142436 6536 142488 6588
rect 160744 6536 160796 6588
rect 174268 6536 174320 6588
rect 345664 6536 345716 6588
rect 138848 6468 138900 6520
rect 159364 6468 159416 6520
rect 186136 6468 186188 6520
rect 371884 6468 371936 6520
rect 148324 6400 148376 6452
rect 434720 6400 434772 6452
rect 155408 6332 155460 6384
rect 466460 6332 466512 6384
rect 144828 6264 144880 6316
rect 173164 6264 173216 6316
rect 219256 6264 219308 6316
rect 572904 6264 572956 6316
rect 147128 6196 147180 6248
rect 518900 6196 518952 6248
rect 101036 6128 101088 6180
rect 181444 6128 181496 6180
rect 187332 6128 187384 6180
rect 572812 6128 572864 6180
rect 81348 5312 81400 5364
rect 128176 5312 128228 5364
rect 69112 5244 69164 5296
rect 96252 5244 96304 5296
rect 96528 5244 96580 5296
rect 193220 5244 193272 5296
rect 232228 5244 232280 5296
rect 412640 5244 412692 5296
rect 86868 5176 86920 5228
rect 285680 5176 285732 5228
rect 31300 5108 31352 5160
rect 270500 5108 270552 5160
rect 68100 5040 68152 5092
rect 214472 5040 214524 5092
rect 235908 5040 235960 5092
rect 481640 5040 481692 5092
rect 68652 4972 68704 5024
rect 171968 4972 172020 5024
rect 177856 4972 177908 5024
rect 207020 4972 207072 5024
rect 207388 4972 207440 5024
rect 455420 4972 455472 5024
rect 65616 4904 65668 4956
rect 137652 4904 137704 4956
rect 143540 4904 143592 4956
rect 550640 4904 550692 4956
rect 572 4836 624 4888
rect 130384 4836 130436 4888
rect 136456 4836 136508 4888
rect 572996 4836 573048 4888
rect 66720 4768 66772 4820
rect 568948 4768 569000 4820
rect 6460 4088 6512 4140
rect 7656 4088 7708 4140
rect 69480 4020 69532 4072
rect 98644 4020 98696 4072
rect 114008 4020 114060 4072
rect 286324 4020 286376 4072
rect 64328 3952 64380 4004
rect 276664 3952 276716 4004
rect 32496 3884 32548 3936
rect 291844 3884 291896 3936
rect 14740 3816 14792 3868
rect 280804 3816 280856 3868
rect 20628 3748 20680 3800
rect 297364 3748 297416 3800
rect 44272 3680 44324 3732
rect 47584 3680 47636 3732
rect 69756 3680 69808 3732
rect 121092 3680 121144 3732
rect 215668 3680 215720 3732
rect 568856 3680 568908 3732
rect 15936 3612 15988 3664
rect 22744 3612 22796 3664
rect 23020 3612 23072 3664
rect 29644 3612 29696 3664
rect 53104 3612 53156 3664
rect 69848 3612 69900 3664
rect 123484 3612 123536 3664
rect 124680 3612 124732 3664
rect 184204 3612 184256 3664
rect 213368 3612 213420 3664
rect 569776 3612 569828 3664
rect 4068 3544 4120 3596
rect 11704 3544 11756 3596
rect 12256 3544 12308 3596
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12348 3476 12400 3528
rect 17040 3544 17092 3596
rect 17868 3544 17920 3596
rect 18236 3544 18288 3596
rect 19248 3544 19300 3596
rect 25320 3544 25372 3596
rect 26148 3544 26200 3596
rect 26884 3544 26936 3596
rect 33600 3544 33652 3596
rect 35164 3544 35216 3596
rect 45468 3544 45520 3596
rect 48964 3544 49016 3596
rect 58624 3544 58676 3596
rect 60832 3544 60884 3596
rect 61936 3544 61988 3596
rect 72424 3544 72476 3596
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 27712 3476 27764 3528
rect 28908 3476 28960 3528
rect 30104 3476 30156 3528
rect 32404 3476 32456 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 38384 3476 38436 3528
rect 39396 3476 39448 3528
rect 39580 3476 39632 3528
rect 40684 3476 40736 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 51356 3476 51408 3528
rect 52368 3476 52420 3528
rect 56048 3476 56100 3528
rect 57152 3476 57204 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 70308 3476 70360 3528
rect 71044 3476 71096 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 73160 3476 73212 3528
rect 73804 3476 73856 3528
rect 95056 3544 95108 3596
rect 89168 3476 89220 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 93952 3476 94004 3528
rect 95148 3476 95200 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 115204 3544 115256 3596
rect 115848 3544 115900 3596
rect 116400 3544 116452 3596
rect 567844 3544 567896 3596
rect 570788 3476 570840 3528
rect 1676 3408 1728 3460
rect 39304 3408 39356 3460
rect 51724 3408 51776 3460
rect 59636 3408 59688 3460
rect 60648 3408 60700 3460
rect 69572 3408 69624 3460
rect 40684 3340 40736 3392
rect 65892 3340 65944 3392
rect 85672 3408 85724 3460
rect 87972 3408 88024 3460
rect 569224 3408 569276 3460
rect 76196 3340 76248 3392
rect 77208 3340 77260 3392
rect 78588 3340 78640 3392
rect 79324 3340 79376 3392
rect 80152 3340 80204 3392
rect 80888 3340 80940 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 102232 3340 102284 3392
rect 122288 3340 122340 3392
rect 122748 3340 122800 3392
rect 125876 3340 125928 3392
rect 126888 3340 126940 3392
rect 126980 3340 127032 3392
rect 128268 3340 128320 3392
rect 149520 3340 149572 3392
rect 150348 3340 150400 3392
rect 151820 3340 151872 3392
rect 153108 3340 153160 3392
rect 184940 3340 184992 3392
rect 186044 3340 186096 3392
rect 189724 3340 189776 3392
rect 190368 3340 190420 3392
rect 196808 3340 196860 3392
rect 197268 3340 197320 3392
rect 199108 3340 199160 3392
rect 200028 3340 200080 3392
rect 206192 3340 206244 3392
rect 206928 3340 206980 3392
rect 218060 3340 218112 3392
rect 219348 3340 219400 3392
rect 223948 3340 224000 3392
rect 224868 3340 224920 3392
rect 225144 3340 225196 3392
rect 226248 3340 226300 3392
rect 229836 3340 229888 3392
rect 230388 3340 230440 3392
rect 234620 3340 234672 3392
rect 235816 3340 235868 3392
rect 28908 3204 28960 3256
rect 33784 3204 33836 3256
rect 2872 3136 2924 3188
rect 4988 3136 5040 3188
rect 7656 3136 7708 3188
rect 10324 3136 10376 3188
rect 19432 3000 19484 3052
rect 21364 3000 21416 3052
rect 47860 3000 47912 3052
rect 50344 3000 50396 3052
rect 52552 3000 52604 3052
rect 54484 3000 54536 3052
rect 69112 2932 69164 2984
rect 71688 2932 71740 2984
rect 24216 2864 24268 2916
rect 24768 2864 24820 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 24320 699718 24348 703520
rect 40512 700330 40540 703520
rect 69848 700460 69900 700466
rect 69848 700402 69900 700408
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 671090 2820 671191
rect 2780 671084 2832 671090
rect 2780 671026 2832 671032
rect 4804 671084 4856 671090
rect 4804 671026 4856 671032
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 2778 580000 2834 580009
rect 2778 579935 2780 579944
rect 2832 579935 2834 579944
rect 2780 579906 2832 579912
rect 3528 576854 3556 619103
rect 3528 576826 3648 576854
rect 3424 567792 3476 567798
rect 3424 567734 3476 567740
rect 3436 514865 3464 567734
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 566370 3556 566879
rect 3620 566506 3648 576826
rect 3608 566500 3660 566506
rect 3608 566442 3660 566448
rect 3516 566364 3568 566370
rect 3516 566306 3568 566312
rect 3514 527912 3570 527921
rect 3514 527847 3570 527856
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 2780 475924 2832 475930
rect 2780 475866 2832 475872
rect 2792 475697 2820 475866
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 2778 423600 2834 423609
rect 2778 423535 2780 423544
rect 2832 423535 2834 423544
rect 2780 423506 2832 423512
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3240 371272 3292 371278
rect 3240 371214 3292 371220
rect 3252 214985 3280 371214
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3238 214976 3294 214985
rect 3238 214911 3294 214920
rect 3344 187746 3372 358391
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 2780 150136 2832 150142
rect 2780 150078 2832 150084
rect 2792 149841 2820 150078
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3332 97980 3384 97986
rect 3332 97922 3384 97928
rect 3344 97617 3372 97922
rect 3330 97608 3386 97617
rect 3330 97543 3386 97552
rect 3436 66570 3464 462567
rect 3528 350538 3556 527847
rect 3976 396092 4028 396098
rect 3976 396034 4028 396040
rect 3700 372632 3752 372638
rect 3700 372574 3752 372580
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3516 350532 3568 350538
rect 3516 350474 3568 350480
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 66842 3556 306167
rect 3620 139398 3648 371311
rect 3712 162897 3740 372574
rect 3884 270564 3936 270570
rect 3884 270506 3936 270512
rect 3790 267200 3846 267209
rect 3790 267135 3846 267144
rect 3698 162888 3754 162897
rect 3698 162823 3754 162832
rect 3608 139392 3660 139398
rect 3608 139334 3660 139340
rect 3606 110664 3662 110673
rect 3606 110599 3662 110608
rect 3516 66836 3568 66842
rect 3516 66778 3568 66784
rect 3424 66564 3476 66570
rect 3424 66506 3476 66512
rect 3620 66230 3648 110599
rect 3804 67318 3832 267135
rect 3896 71641 3924 270506
rect 3988 201929 4016 396034
rect 4066 254144 4122 254153
rect 4066 254079 4122 254088
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3882 71632 3938 71641
rect 3882 71567 3938 71576
rect 4080 67454 4108 254079
rect 4816 67522 4844 671026
rect 4896 579964 4948 579970
rect 4896 579906 4948 579912
rect 4908 67590 4936 579906
rect 10324 570988 10376 570994
rect 10324 570930 10376 570936
rect 5080 568064 5132 568070
rect 5080 568006 5132 568012
rect 4988 560312 5040 560318
rect 4988 560254 5040 560260
rect 5000 150142 5028 560254
rect 5092 475930 5120 568006
rect 7656 567996 7708 568002
rect 7656 567938 7708 567944
rect 7564 566364 7616 566370
rect 7564 566306 7616 566312
rect 5080 475924 5132 475930
rect 5080 475866 5132 475872
rect 5080 423564 5132 423570
rect 5080 423506 5132 423512
rect 4988 150136 5040 150142
rect 4988 150078 5040 150084
rect 4988 69692 5040 69698
rect 4988 69634 5040 69640
rect 4896 67584 4948 67590
rect 4896 67526 4948 67532
rect 4804 67516 4856 67522
rect 4804 67458 4856 67464
rect 4068 67448 4120 67454
rect 4068 67390 4120 67396
rect 3792 67312 3844 67318
rect 3792 67254 3844 67260
rect 3700 66904 3752 66910
rect 3700 66846 3752 66852
rect 3608 66224 3660 66230
rect 3608 66166 3660 66172
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3712 32473 3740 66846
rect 3698 32464 3754 32473
rect 3698 32399 3754 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2884 480 2912 3130
rect 4080 480 4108 3538
rect 5000 3194 5028 69634
rect 5092 67250 5120 423506
rect 5540 396772 5592 396778
rect 5540 396714 5592 396720
rect 5552 393314 5580 396714
rect 5184 393286 5580 393314
rect 5184 371278 5212 393286
rect 5172 371272 5224 371278
rect 5172 371214 5224 371220
rect 5172 187740 5224 187746
rect 5172 187682 5224 187688
rect 5184 175250 5212 187682
rect 5184 175222 5580 175250
rect 5552 171154 5580 175222
rect 5540 171148 5592 171154
rect 5540 171090 5592 171096
rect 7576 67386 7604 566306
rect 7668 320142 7696 567938
rect 7656 320136 7708 320142
rect 7656 320078 7708 320084
rect 9588 176724 9640 176730
rect 9588 176666 9640 176672
rect 8300 171080 8352 171086
rect 8300 171022 8352 171028
rect 8312 168434 8340 171022
rect 8300 168428 8352 168434
rect 8300 168370 8352 168376
rect 7656 69760 7708 69766
rect 7656 69702 7708 69708
rect 7564 67380 7616 67386
rect 7564 67322 7616 67328
rect 5080 67244 5132 67250
rect 5080 67186 5132 67192
rect 7668 4146 7696 69702
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 6472 480 6500 4082
rect 9600 3534 9628 176666
rect 9772 168428 9824 168434
rect 9772 168370 9824 168376
rect 9784 164286 9812 168370
rect 9772 164280 9824 164286
rect 9772 164222 9824 164228
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7668 480 7696 3130
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 10336 3194 10364 570930
rect 12348 570648 12400 570654
rect 12348 570590 12400 570596
rect 11704 568200 11756 568206
rect 11704 568142 11756 568148
rect 10416 568132 10468 568138
rect 10416 568074 10468 568080
rect 10428 97986 10456 568074
rect 10968 231872 11020 231878
rect 10968 231814 11020 231820
rect 10416 97980 10468 97986
rect 10416 97922 10468 97928
rect 10980 3534 11008 231814
rect 11716 3602 11744 568142
rect 11796 567656 11848 567662
rect 11796 567598 11848 567604
rect 11808 59362 11836 567598
rect 11796 59356 11848 59362
rect 11796 59298 11848 59304
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 11164 480 11192 3470
rect 12268 1850 12296 3538
rect 12360 3534 12388 570590
rect 22744 570444 22796 570450
rect 22744 570386 22796 570392
rect 21364 417376 21416 417382
rect 21364 417318 21416 417324
rect 13728 411324 13780 411330
rect 13728 411266 13780 411272
rect 12440 400240 12492 400246
rect 12440 400182 12492 400188
rect 12452 396778 12480 400182
rect 12440 396772 12492 396778
rect 12440 396714 12492 396720
rect 13740 6914 13768 411266
rect 21376 408814 21404 417318
rect 18604 408808 18656 408814
rect 18604 408750 18656 408756
rect 21364 408808 21416 408814
rect 21364 408750 21416 408756
rect 18616 407250 18644 408750
rect 15844 407244 15896 407250
rect 15844 407186 15896 407192
rect 18604 407244 18656 407250
rect 18604 407186 18656 407192
rect 15856 400246 15884 407186
rect 15844 400240 15896 400246
rect 15844 400182 15896 400188
rect 15200 164212 15252 164218
rect 15200 164154 15252 164160
rect 15212 161430 15240 164154
rect 15200 161424 15252 161430
rect 15200 161366 15252 161372
rect 19248 161424 19300 161430
rect 19248 161366 19300 161372
rect 19260 154442 19288 161366
rect 19260 154414 19380 154442
rect 19352 151842 19380 154414
rect 19340 151836 19392 151842
rect 19340 151778 19392 151784
rect 22008 98048 22060 98054
rect 22008 97990 22060 97996
rect 21364 69828 21416 69834
rect 21364 69770 21416 69776
rect 19248 65952 19300 65958
rect 19248 65894 19300 65900
rect 17868 65272 17920 65278
rect 17868 65214 17920 65220
rect 13556 6886 13768 6914
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14740 3868 14792 3874
rect 14740 3810 14792 3816
rect 14752 480 14780 3810
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15948 480 15976 3606
rect 17880 3602 17908 65214
rect 19260 3602 19288 65894
rect 20628 3800 20680 3806
rect 20628 3742 20680 3748
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 17052 480 17080 3538
rect 18248 480 18276 3538
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 20640 480 20668 3742
rect 21376 3058 21404 69770
rect 22020 6914 22048 97990
rect 21836 6886 22048 6914
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21836 480 21864 6886
rect 22756 3670 22784 570386
rect 24124 466472 24176 466478
rect 24124 466414 24176 466420
rect 24136 424794 24164 466414
rect 22836 424788 22888 424794
rect 22836 424730 22888 424736
rect 24124 424788 24176 424794
rect 24124 424730 24176 424736
rect 22848 417382 22876 424730
rect 22836 417376 22888 417382
rect 22836 417318 22888 417324
rect 24780 327078 24808 699654
rect 68744 630692 68796 630698
rect 68744 630634 68796 630640
rect 64144 571056 64196 571062
rect 64144 570998 64196 571004
rect 58624 570852 58676 570858
rect 58624 570794 58676 570800
rect 57244 570784 57296 570790
rect 57244 570726 57296 570732
rect 54484 570716 54536 570722
rect 54484 570658 54536 570664
rect 39304 570308 39356 570314
rect 39304 570250 39356 570256
rect 26884 570036 26936 570042
rect 26884 569978 26936 569984
rect 25136 469872 25188 469878
rect 25136 469814 25188 469820
rect 25148 466478 25176 469814
rect 25136 466472 25188 466478
rect 25136 466414 25188 466420
rect 24768 327072 24820 327078
rect 24768 327014 24820 327020
rect 26148 208412 26200 208418
rect 26148 208354 26200 208360
rect 22836 151768 22888 151774
rect 22836 151710 22888 151716
rect 22848 138718 22876 151710
rect 22836 138712 22888 138718
rect 22836 138654 22888 138660
rect 24124 138712 24176 138718
rect 24124 138654 24176 138660
rect 24136 129810 24164 138654
rect 24124 129804 24176 129810
rect 24124 129746 24176 129752
rect 24768 65884 24820 65890
rect 24768 65826 24820 65832
rect 22744 3664 22796 3670
rect 22744 3606 22796 3612
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 23032 480 23060 3606
rect 24780 2922 24808 65826
rect 26160 3602 26188 208354
rect 26896 3602 26924 569978
rect 37188 510604 37240 510610
rect 37188 510546 37240 510552
rect 37200 502994 37228 510546
rect 35164 502988 35216 502994
rect 35164 502930 35216 502936
rect 37188 502988 37240 502994
rect 37188 502930 37240 502936
rect 35176 491298 35204 502930
rect 33232 491292 33284 491298
rect 33232 491234 33284 491240
rect 35164 491292 35216 491298
rect 35164 491234 35216 491240
rect 33244 487218 33272 491234
rect 32404 487212 32456 487218
rect 32404 487154 32456 487160
rect 33232 487212 33284 487218
rect 33232 487154 33284 487160
rect 32416 478922 32444 487154
rect 30380 478916 30432 478922
rect 30380 478858 30432 478864
rect 32404 478916 32456 478922
rect 32404 478858 32456 478864
rect 30392 470594 30420 478858
rect 30024 470566 30420 470594
rect 30024 469878 30052 470566
rect 30012 469872 30064 469878
rect 30012 469814 30064 469820
rect 27528 302932 27580 302938
rect 27528 302874 27580 302880
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 24216 2916 24268 2922
rect 24216 2858 24268 2864
rect 24768 2916 24820 2922
rect 24768 2858 24820 2864
rect 24228 480 24256 2858
rect 25332 480 25360 3538
rect 27540 3534 27568 302874
rect 28264 129736 28316 129742
rect 28264 129678 28316 129684
rect 28276 125594 28304 129678
rect 28264 125588 28316 125594
rect 28264 125530 28316 125536
rect 30288 125588 30340 125594
rect 30288 125530 30340 125536
rect 30300 122834 30328 125530
rect 30300 122806 30420 122834
rect 30392 118182 30420 122806
rect 30380 118176 30432 118182
rect 30380 118118 30432 118124
rect 32404 118176 32456 118182
rect 32404 118118 32456 118124
rect 32416 105534 32444 118118
rect 32404 105528 32456 105534
rect 32404 105470 32456 105476
rect 37280 105528 37332 105534
rect 37280 105470 37332 105476
rect 37292 100910 37320 105470
rect 37280 100904 37332 100910
rect 37280 100846 37332 100852
rect 37188 82884 37240 82890
rect 37188 82826 37240 82832
rect 37096 69964 37148 69970
rect 37096 69906 37148 69912
rect 35808 69896 35860 69902
rect 35808 69838 35860 69844
rect 32404 66156 32456 66162
rect 32404 66098 32456 66104
rect 29644 65612 29696 65618
rect 29644 65554 29696 65560
rect 28908 65340 28960 65346
rect 28908 65282 28960 65288
rect 28920 3534 28948 65282
rect 29656 3670 29684 65554
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 26528 480 26556 3470
rect 27724 480 27752 3470
rect 28908 3256 28960 3262
rect 28908 3198 28960 3204
rect 28920 480 28948 3198
rect 30116 480 30144 3470
rect 31312 480 31340 5102
rect 32416 3534 32444 66098
rect 33784 65204 33836 65210
rect 33784 65146 33836 65152
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 32508 1986 32536 3878
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 32416 1958 32536 1986
rect 32416 480 32444 1958
rect 33612 480 33640 3538
rect 33796 3262 33824 65146
rect 35164 65136 35216 65142
rect 35164 65078 35216 65084
rect 35176 3602 35204 65078
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 35820 3534 35848 69838
rect 37108 3534 37136 69906
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 33784 3256 33836 3262
rect 33784 3198 33836 3204
rect 34808 480 34836 3470
rect 36004 480 36032 3470
rect 37200 480 37228 82826
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 38396 480 38424 3470
rect 39316 3466 39344 570250
rect 50344 570240 50396 570246
rect 50344 570182 50396 570188
rect 46848 567860 46900 567866
rect 46848 567802 46900 567808
rect 44088 567724 44140 567730
rect 44088 567666 44140 567672
rect 39396 567384 39448 567390
rect 39396 567326 39448 567332
rect 39408 3534 39436 567326
rect 42064 532092 42116 532098
rect 42064 532034 42116 532040
rect 42076 514826 42104 532034
rect 39672 514820 39724 514826
rect 39672 514762 39724 514768
rect 42064 514820 42116 514826
rect 42064 514762 42116 514768
rect 39684 510678 39712 514762
rect 39672 510672 39724 510678
rect 39672 510614 39724 510620
rect 40040 100904 40092 100910
rect 40040 100846 40092 100852
rect 40052 95198 40080 100846
rect 40040 95192 40092 95198
rect 40040 95134 40092 95140
rect 42616 95192 42668 95198
rect 42616 95134 42668 95140
rect 42628 92342 42656 95134
rect 42616 92336 42668 92342
rect 42616 92278 42668 92284
rect 42708 70032 42760 70038
rect 42708 69974 42760 69980
rect 40684 65476 40736 65482
rect 40684 65418 40736 65424
rect 40696 3534 40724 65418
rect 42720 3534 42748 69974
rect 44100 3534 44128 567666
rect 44180 92336 44232 92342
rect 44180 92278 44232 92284
rect 44192 90370 44220 92278
rect 44180 90364 44232 90370
rect 44180 90306 44232 90312
rect 46860 6914 46888 567802
rect 47584 546440 47636 546446
rect 47584 546382 47636 546388
rect 47596 532098 47624 546382
rect 47584 532092 47636 532098
rect 47584 532034 47636 532040
rect 49608 90364 49660 90370
rect 49608 90306 49660 90312
rect 49620 89706 49648 90306
rect 49620 89678 49740 89706
rect 49712 86970 49740 89678
rect 49700 86964 49752 86970
rect 49700 86906 49752 86912
rect 47584 65544 47636 65550
rect 47584 65486 47636 65492
rect 46676 6886 46888 6914
rect 44272 3732 44324 3738
rect 44272 3674 44324 3680
rect 39396 3528 39448 3534
rect 39396 3470 39448 3476
rect 39580 3528 39632 3534
rect 39580 3470 39632 3476
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 39304 3460 39356 3466
rect 39304 3402 39356 3408
rect 39592 480 39620 3470
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3674
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45480 480 45508 3538
rect 46676 480 46704 6886
rect 47596 3738 47624 65486
rect 47584 3732 47636 3738
rect 47584 3674 47636 3680
rect 48964 3596 49016 3602
rect 48964 3538 49016 3544
rect 47860 3052 47912 3058
rect 47860 2994 47912 3000
rect 47872 480 47900 2994
rect 48976 480 49004 3538
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50172 480 50200 3470
rect 50356 3058 50384 570182
rect 50436 409896 50488 409902
rect 50436 409838 50488 409844
rect 50448 66026 50476 409838
rect 52368 342916 52420 342922
rect 52368 342858 52420 342864
rect 52276 86964 52328 86970
rect 52276 86906 52328 86912
rect 52288 82482 52316 86906
rect 52276 82476 52328 82482
rect 52276 82418 52328 82424
rect 50988 70100 51040 70106
rect 50988 70042 51040 70048
rect 50436 66020 50488 66026
rect 50436 65962 50488 65968
rect 51000 3534 51028 70042
rect 51724 65816 51776 65822
rect 51724 65758 51776 65764
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 50344 3052 50396 3058
rect 50344 2994 50396 3000
rect 51368 480 51396 3470
rect 51736 3466 51764 65758
rect 52380 3534 52408 342858
rect 53748 66088 53800 66094
rect 53748 66030 53800 66036
rect 53104 65680 53156 65686
rect 53104 65622 53156 65628
rect 53116 3670 53144 65622
rect 53104 3664 53156 3670
rect 53104 3606 53156 3612
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 51724 3460 51776 3466
rect 51724 3402 51776 3408
rect 52552 3052 52604 3058
rect 52552 2994 52604 3000
rect 52564 480 52592 2994
rect 53760 480 53788 66030
rect 54496 3058 54524 570658
rect 55864 551812 55916 551818
rect 55864 551754 55916 551760
rect 55876 546514 55904 551754
rect 55864 546508 55916 546514
rect 55864 546450 55916 546456
rect 55128 364404 55180 364410
rect 55128 364346 55180 364352
rect 55140 6914 55168 364346
rect 56508 82476 56560 82482
rect 56508 82418 56560 82424
rect 56520 77314 56548 82418
rect 56508 77308 56560 77314
rect 56508 77250 56560 77256
rect 57256 6914 57284 570726
rect 57888 556232 57940 556238
rect 57888 556174 57940 556180
rect 57900 551818 57928 556174
rect 57888 551812 57940 551818
rect 57888 551754 57940 551760
rect 57888 69624 57940 69630
rect 57888 69566 57940 69572
rect 54956 6886 55168 6914
rect 57164 6886 57284 6914
rect 54484 3052 54536 3058
rect 54484 2994 54536 3000
rect 54956 480 54984 6886
rect 57164 3534 57192 6886
rect 57900 3534 57928 69566
rect 58636 3602 58664 570794
rect 62028 567588 62080 567594
rect 62028 567530 62080 567536
rect 61936 69420 61988 69426
rect 61936 69362 61988 69368
rect 60648 65748 60700 65754
rect 60648 65690 60700 65696
rect 59268 44192 59320 44198
rect 59268 44134 59320 44140
rect 58624 3596 58676 3602
rect 58624 3538 58676 3544
rect 59280 3534 59308 44134
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 57152 3528 57204 3534
rect 57152 3470 57204 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 60660 3466 60688 65690
rect 61948 16574 61976 69362
rect 61856 16546 61976 16574
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 59636 3460 59688 3466
rect 59636 3402 59688 3408
rect 60648 3460 60700 3466
rect 60648 3402 60700 3408
rect 59648 480 59676 3402
rect 60844 480 60872 3538
rect 61856 3482 61884 16546
rect 62040 6914 62068 567530
rect 63408 238808 63460 238814
rect 63408 238750 63460 238756
rect 63420 6914 63448 238750
rect 63500 77240 63552 77246
rect 63500 77182 63552 77188
rect 63512 75206 63540 77182
rect 63500 75200 63552 75206
rect 63500 75142 63552 75148
rect 64156 44198 64184 570998
rect 65524 570580 65576 570586
rect 65524 570522 65576 570528
rect 64880 559904 64932 559910
rect 64880 559846 64932 559852
rect 64892 557546 64920 559846
rect 64800 557518 64920 557546
rect 64800 556238 64828 557518
rect 64788 556232 64840 556238
rect 64788 556174 64840 556180
rect 65536 342922 65564 570522
rect 66076 570104 66128 570110
rect 66076 570046 66128 570052
rect 65984 536852 66036 536858
rect 65984 536794 66036 536800
rect 65800 426488 65852 426494
rect 65800 426430 65852 426436
rect 65708 356108 65760 356114
rect 65708 356050 65760 356056
rect 65524 342916 65576 342922
rect 65524 342858 65576 342864
rect 65524 302252 65576 302258
rect 65524 302194 65576 302200
rect 65432 161560 65484 161566
rect 65432 161502 65484 161508
rect 65340 69352 65392 69358
rect 65340 69294 65392 69300
rect 64144 44192 64196 44198
rect 64144 44134 64196 44140
rect 65352 16574 65380 69294
rect 65444 67862 65472 161502
rect 65432 67856 65484 67862
rect 65432 67798 65484 67804
rect 65536 62830 65564 302194
rect 65616 285728 65668 285734
rect 65616 285670 65668 285676
rect 65524 62824 65576 62830
rect 65524 62766 65576 62772
rect 65352 16546 65564 16574
rect 61948 6886 62068 6914
rect 63236 6886 63448 6914
rect 61948 3602 61976 6886
rect 61936 3596 61988 3602
rect 61936 3538 61988 3544
rect 61856 3454 62068 3482
rect 62040 480 62068 3454
rect 63236 480 63264 6886
rect 64328 4004 64380 4010
rect 64328 3946 64380 3952
rect 64340 480 64368 3946
rect 65536 480 65564 16546
rect 65628 4962 65656 285670
rect 65720 68338 65748 356050
rect 65708 68332 65760 68338
rect 65708 68274 65760 68280
rect 65812 67930 65840 426430
rect 65892 403300 65944 403306
rect 65892 403242 65944 403248
rect 65800 67924 65852 67930
rect 65800 67866 65852 67872
rect 65616 4956 65668 4962
rect 65616 4898 65668 4904
rect 65904 3398 65932 403242
rect 65996 67046 66024 536794
rect 66088 68406 66116 570046
rect 66168 567316 66220 567322
rect 66168 567258 66220 567264
rect 66076 68400 66128 68406
rect 66076 68342 66128 68348
rect 65984 67040 66036 67046
rect 65984 66982 66036 66988
rect 66180 66706 66208 567258
rect 68652 561740 68704 561746
rect 68652 561682 68704 561688
rect 67638 560416 67694 560425
rect 67638 560351 67694 560360
rect 67652 560318 67680 560351
rect 67640 560312 67692 560318
rect 67640 560254 67692 560260
rect 68664 559910 68692 561682
rect 68652 559904 68704 559910
rect 68652 559846 68704 559852
rect 68756 552537 68784 630634
rect 68836 570512 68888 570518
rect 68836 570454 68888 570460
rect 68742 552528 68798 552537
rect 68742 552463 68798 552472
rect 67546 544912 67602 544921
rect 67546 544847 67602 544856
rect 67454 529136 67510 529145
rect 67454 529071 67510 529080
rect 67362 521248 67418 521257
rect 67362 521183 67418 521192
rect 67270 505744 67326 505753
rect 67270 505679 67326 505688
rect 67178 435296 67234 435305
rect 67178 435231 67234 435240
rect 67086 419792 67142 419801
rect 67086 419727 67142 419736
rect 66994 224224 67050 224233
rect 66994 224159 67050 224168
rect 66902 185328 66958 185337
rect 66902 185263 66958 185272
rect 66812 129804 66864 129810
rect 66812 129746 66864 129752
rect 66824 68542 66852 129746
rect 66812 68536 66864 68542
rect 66812 68478 66864 68484
rect 66916 68270 66944 185263
rect 67008 68746 67036 224159
rect 66996 68740 67048 68746
rect 66996 68682 67048 68688
rect 66904 68264 66956 68270
rect 66904 68206 66956 68212
rect 67100 66978 67128 419727
rect 67192 68202 67220 435231
rect 67180 68196 67232 68202
rect 67180 68138 67232 68144
rect 67284 67794 67312 505679
rect 67376 68134 67404 521183
rect 67364 68128 67416 68134
rect 67364 68070 67416 68076
rect 67272 67788 67324 67794
rect 67272 67730 67324 67736
rect 67088 66972 67140 66978
rect 67088 66914 67140 66920
rect 67468 66774 67496 529071
rect 67456 66768 67508 66774
rect 67456 66710 67508 66716
rect 66168 66700 66220 66706
rect 66168 66642 66220 66648
rect 67560 55894 67588 544847
rect 67638 537024 67694 537033
rect 67638 536959 67694 536968
rect 67652 536858 67680 536959
rect 67640 536852 67692 536858
rect 67640 536794 67692 536800
rect 68742 513632 68798 513641
rect 68742 513567 68798 513576
rect 68650 497856 68706 497865
rect 68650 497791 68706 497800
rect 68374 482352 68430 482361
rect 68374 482287 68430 482296
rect 68282 474464 68338 474473
rect 68282 474399 68338 474408
rect 67914 427408 67970 427417
rect 67914 427343 67970 427352
rect 67928 426494 67956 427343
rect 67916 426488 67968 426494
rect 67916 426430 67968 426436
rect 67638 411904 67694 411913
rect 67638 411839 67694 411848
rect 67652 411330 67680 411839
rect 67640 411324 67692 411330
rect 67640 411266 67692 411272
rect 68006 404016 68062 404025
rect 68006 403951 68062 403960
rect 68020 403306 68048 403951
rect 68008 403300 68060 403306
rect 68008 403242 68060 403248
rect 67638 396400 67694 396409
rect 67638 396335 67694 396344
rect 67652 396098 67680 396335
rect 67640 396092 67692 396098
rect 67640 396034 67692 396040
rect 67638 372736 67694 372745
rect 67638 372671 67694 372680
rect 67652 372638 67680 372671
rect 67640 372632 67692 372638
rect 67640 372574 67692 372580
rect 67638 365120 67694 365129
rect 67638 365055 67694 365064
rect 67652 364410 67680 365055
rect 67640 364404 67692 364410
rect 67640 364346 67692 364352
rect 67822 357232 67878 357241
rect 67822 357167 67878 357176
rect 67836 356114 67864 357167
rect 67824 356108 67876 356114
rect 67824 356050 67876 356056
rect 67640 350532 67692 350538
rect 67640 350474 67692 350480
rect 67652 349353 67680 350474
rect 67638 349344 67694 349353
rect 67638 349279 67694 349288
rect 67640 327072 67692 327078
rect 67640 327014 67692 327020
rect 67652 325961 67680 327014
rect 67638 325952 67694 325961
rect 67638 325887 67694 325896
rect 68192 310480 68244 310486
rect 68192 310422 68244 310428
rect 67822 302560 67878 302569
rect 67822 302495 67878 302504
rect 67836 302258 67864 302495
rect 67824 302252 67876 302258
rect 67824 302194 67876 302200
rect 67822 286784 67878 286793
rect 67822 286719 67878 286728
rect 67836 285734 67864 286719
rect 67824 285728 67876 285734
rect 67824 285670 67876 285676
rect 68204 278905 68232 310422
rect 68296 302938 68324 474399
rect 68284 302932 68336 302938
rect 68284 302874 68336 302880
rect 68190 278896 68246 278905
rect 68190 278831 68246 278840
rect 67638 271280 67694 271289
rect 67638 271215 67694 271224
rect 67652 270570 67680 271215
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 68282 263392 68338 263401
rect 68282 263327 68338 263336
rect 68190 255504 68246 255513
rect 68190 255439 68246 255448
rect 67638 240000 67694 240009
rect 67638 239935 67694 239944
rect 67652 238814 67680 239935
rect 67640 238808 67692 238814
rect 67640 238750 67692 238756
rect 67638 232112 67694 232121
rect 67638 232047 67694 232056
rect 67652 231878 67680 232047
rect 67640 231872 67692 231878
rect 67640 231814 67692 231820
rect 67638 208720 67694 208729
rect 67638 208655 67694 208664
rect 67652 208418 67680 208655
rect 67640 208412 67692 208418
rect 67640 208354 67692 208360
rect 67730 200832 67786 200841
rect 67730 200767 67786 200776
rect 67638 177440 67694 177449
rect 67638 177375 67694 177384
rect 67652 176730 67680 177375
rect 67640 176724 67692 176730
rect 67640 176666 67692 176672
rect 67638 161664 67694 161673
rect 67638 161599 67694 161608
rect 67652 161566 67680 161599
rect 67640 161560 67692 161566
rect 67640 161502 67692 161508
rect 67640 139392 67692 139398
rect 67640 139334 67692 139340
rect 67652 138281 67680 139334
rect 67638 138272 67694 138281
rect 67638 138207 67694 138216
rect 67638 130384 67694 130393
rect 67638 130319 67694 130328
rect 67652 129810 67680 130319
rect 67640 129804 67692 129810
rect 67640 129746 67692 129752
rect 67638 99104 67694 99113
rect 67638 99039 67694 99048
rect 67652 98054 67680 99039
rect 67640 98048 67692 98054
rect 67640 97990 67692 97996
rect 67638 91488 67694 91497
rect 67638 91423 67694 91432
rect 67652 69494 67680 91423
rect 67640 69488 67692 69494
rect 67640 69430 67692 69436
rect 67744 68950 67772 200767
rect 68098 192944 68154 192953
rect 68098 192879 68154 192888
rect 68006 154048 68062 154057
rect 68006 153983 68062 153992
rect 67914 146160 67970 146169
rect 67914 146095 67970 146104
rect 67822 114880 67878 114889
rect 67822 114815 67878 114824
rect 67732 68944 67784 68950
rect 67732 68886 67784 68892
rect 67836 68610 67864 114815
rect 67928 68882 67956 146095
rect 67916 68876 67968 68882
rect 67916 68818 67968 68824
rect 67824 68604 67876 68610
rect 67824 68546 67876 68552
rect 68020 67726 68048 153983
rect 68112 146266 68140 192879
rect 68100 146260 68152 146266
rect 68100 146202 68152 146208
rect 68098 122768 68154 122777
rect 68098 122703 68154 122712
rect 68008 67720 68060 67726
rect 68008 67662 68060 67668
rect 67548 55888 67600 55894
rect 67548 55830 67600 55836
rect 68112 5098 68140 122703
rect 68204 66638 68232 255439
rect 68192 66632 68244 66638
rect 68192 66574 68244 66580
rect 68296 57254 68324 263327
rect 68388 247722 68416 482287
rect 68558 466576 68614 466585
rect 68558 466511 68614 466520
rect 68466 443184 68522 443193
rect 68466 443119 68522 443128
rect 68376 247716 68428 247722
rect 68376 247658 68428 247664
rect 68374 247616 68430 247625
rect 68374 247551 68430 247560
rect 68388 193186 68416 247551
rect 68376 193180 68428 193186
rect 68376 193122 68428 193128
rect 68374 83600 68430 83609
rect 68374 83535 68430 83544
rect 68388 82890 68416 83535
rect 68376 82884 68428 82890
rect 68376 82826 68428 82832
rect 68376 69012 68428 69018
rect 68376 68954 68428 68960
rect 68388 67658 68416 68954
rect 68376 67652 68428 67658
rect 68376 67594 68428 67600
rect 68480 64394 68508 443119
rect 68572 68678 68600 466511
rect 68664 451178 68692 497791
rect 68652 451172 68704 451178
rect 68652 451114 68704 451120
rect 68650 451072 68706 451081
rect 68650 451007 68706 451016
rect 68560 68672 68612 68678
rect 68560 68614 68612 68620
rect 68468 64388 68520 64394
rect 68468 64330 68520 64336
rect 68284 57248 68336 57254
rect 68284 57190 68336 57196
rect 68100 5092 68152 5098
rect 68100 5034 68152 5040
rect 68664 5030 68692 451007
rect 68756 69154 68784 513567
rect 68744 69148 68796 69154
rect 68744 69090 68796 69096
rect 68744 69012 68796 69018
rect 68744 68954 68796 68960
rect 68756 68066 68784 68954
rect 68848 68474 68876 570454
rect 69664 570172 69716 570178
rect 69664 570114 69716 570120
rect 68928 569968 68980 569974
rect 68928 569910 68980 569916
rect 68940 69018 68968 569910
rect 69020 565888 69072 565894
rect 69020 565830 69072 565836
rect 69032 561746 69060 565830
rect 69020 561740 69072 561746
rect 69020 561682 69072 561688
rect 69018 388512 69074 388521
rect 69018 388447 69074 388456
rect 69032 69562 69060 388447
rect 69202 318064 69258 318073
rect 69202 317999 69258 318008
rect 69110 310176 69166 310185
rect 69110 310111 69166 310120
rect 69020 69556 69072 69562
rect 69020 69498 69072 69504
rect 68928 69012 68980 69018
rect 68928 68954 68980 68960
rect 68928 68808 68980 68814
rect 68928 68750 68980 68756
rect 68836 68468 68888 68474
rect 68836 68410 68888 68416
rect 68744 68060 68796 68066
rect 68744 68002 68796 68008
rect 68652 5024 68704 5030
rect 68652 4966 68704 4972
rect 66720 4820 66772 4826
rect 66720 4762 66772 4768
rect 65892 3392 65944 3398
rect 65892 3334 65944 3340
rect 66732 480 66760 4762
rect 68940 3534 68968 68750
rect 69124 5302 69152 310111
rect 69216 67998 69244 317999
rect 69294 294672 69350 294681
rect 69294 294607 69350 294616
rect 69308 68746 69336 294607
rect 69572 193180 69624 193186
rect 69572 193122 69624 193128
rect 69480 146260 69532 146266
rect 69480 146202 69532 146208
rect 69388 75200 69440 75206
rect 69388 75142 69440 75148
rect 69400 69290 69428 75142
rect 69388 69284 69440 69290
rect 69388 69226 69440 69232
rect 69296 68740 69348 68746
rect 69296 68682 69348 68688
rect 69204 67992 69256 67998
rect 69204 67934 69256 67940
rect 69112 5296 69164 5302
rect 69112 5238 69164 5244
rect 69492 4078 69520 146202
rect 69480 4072 69532 4078
rect 69480 4014 69532 4020
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 67928 480 67956 3470
rect 69584 3466 69612 193122
rect 69676 68814 69704 570114
rect 69756 451172 69808 451178
rect 69756 451114 69808 451120
rect 69664 68808 69716 68814
rect 69664 68750 69716 68756
rect 69768 3738 69796 451114
rect 69860 310486 69888 700402
rect 89180 700398 89208 703520
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 105464 699825 105492 703520
rect 154132 700670 154160 703520
rect 170324 700738 170352 703520
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 218992 700330 219020 703520
rect 105544 700324 105596 700330
rect 105544 700266 105596 700272
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 105450 699816 105506 699825
rect 105450 699751 105506 699760
rect 105556 571334 105584 700266
rect 235184 699825 235212 703520
rect 283852 700874 283880 703520
rect 283840 700868 283892 700874
rect 283840 700810 283892 700816
rect 300136 700602 300164 703520
rect 318708 700800 318760 700806
rect 318708 700742 318760 700748
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 277308 700528 277360 700534
rect 277308 700470 277360 700476
rect 235170 699816 235226 699825
rect 235170 699751 235226 699760
rect 256608 616888 256660 616894
rect 256608 616830 256660 616836
rect 105544 571328 105596 571334
rect 105544 571270 105596 571276
rect 107200 571328 107252 571334
rect 107200 571270 107252 571276
rect 249982 571296 250038 571305
rect 75368 569968 75420 569974
rect 75368 569910 75420 569916
rect 75380 567868 75408 569910
rect 107212 567868 107240 571270
rect 249982 571231 250038 571240
rect 186504 571056 186556 571062
rect 176014 571024 176070 571033
rect 186504 570998 186556 571004
rect 176014 570959 176070 570968
rect 138848 570852 138900 570858
rect 138848 570794 138900 570800
rect 123024 570648 123076 570654
rect 123024 570590 123076 570596
rect 123036 567868 123064 570590
rect 138860 567868 138888 570794
rect 149520 570784 149572 570790
rect 149520 570726 149572 570732
rect 149532 567868 149560 570726
rect 165344 570716 165396 570722
rect 165344 570658 165396 570664
rect 165356 567868 165384 570658
rect 176028 567868 176056 570959
rect 178132 570376 178184 570382
rect 178132 570318 178184 570324
rect 178144 568585 178172 570318
rect 178130 568576 178186 568585
rect 178130 568511 178186 568520
rect 186516 567868 186544 570998
rect 191840 570580 191892 570586
rect 191840 570522 191892 570528
rect 191852 567868 191880 570522
rect 239312 570512 239364 570518
rect 239312 570454 239364 570460
rect 196992 570444 197044 570450
rect 196992 570386 197044 570392
rect 197004 567868 197032 570386
rect 234160 568268 234212 568274
rect 234160 568210 234212 568216
rect 218336 568064 218388 568070
rect 218336 568006 218388 568012
rect 223304 568064 223356 568070
rect 223304 568006 223356 568012
rect 208032 567928 208084 567934
rect 207690 567876 208032 567882
rect 218348 567882 218376 568006
rect 207690 567870 208084 567876
rect 207690 567854 208072 567870
rect 218178 567854 218376 567882
rect 223316 567882 223344 568006
rect 223316 567854 223514 567882
rect 234172 567868 234200 568210
rect 239324 567868 239352 570454
rect 249996 567868 250024 571231
rect 256620 570790 256648 616830
rect 277320 571334 277348 700470
rect 276480 571328 276532 571334
rect 276480 571270 276532 571276
rect 277308 571328 277360 571334
rect 277308 571270 277360 571276
rect 255320 570784 255372 570790
rect 255320 570726 255372 570732
rect 256608 570784 256660 570790
rect 256608 570726 256660 570732
rect 255332 567868 255360 570726
rect 276492 567868 276520 571270
rect 302790 571160 302846 571169
rect 302790 571095 302846 571104
rect 292302 570888 292358 570897
rect 292302 570823 292358 570832
rect 286966 570752 287022 570761
rect 286966 570687 287022 570696
rect 286980 567868 287008 570687
rect 292316 567868 292344 570823
rect 297454 570616 297510 570625
rect 297454 570551 297510 570560
rect 297468 567868 297496 570551
rect 302804 567868 302832 571095
rect 318720 567882 318748 700742
rect 348804 700738 348832 703520
rect 333980 700732 334032 700738
rect 333980 700674 334032 700680
rect 348792 700732 348844 700738
rect 348792 700674 348844 700680
rect 333992 576854 334020 700674
rect 364996 700466 365024 703520
rect 413664 700466 413692 703520
rect 418160 700664 418212 700670
rect 418160 700606 418212 700612
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 418172 576854 418200 700606
rect 424324 700392 424376 700398
rect 424324 700334 424376 700340
rect 333992 576826 334296 576854
rect 418172 576826 418752 576854
rect 318642 567854 318748 567882
rect 334268 567882 334296 576826
rect 392766 571024 392822 571033
rect 392766 570959 392822 570968
rect 349986 570888 350042 570897
rect 349986 570823 350042 570832
rect 350000 570625 350028 570823
rect 376942 570752 376998 570761
rect 376942 570687 376998 570696
rect 349986 570616 350042 570625
rect 349986 570551 350042 570560
rect 350448 570308 350500 570314
rect 350448 570250 350500 570256
rect 334268 567854 334650 567882
rect 350460 567868 350488 570250
rect 355784 568200 355836 568206
rect 355784 568142 355836 568148
rect 355796 567868 355824 568142
rect 360936 568132 360988 568138
rect 360936 568074 360988 568080
rect 360948 567868 360976 568074
rect 365996 567996 366048 568002
rect 365996 567938 366048 567944
rect 371976 567996 372028 568002
rect 371976 567938 372028 567944
rect 366008 567882 366036 567938
rect 371988 567882 372016 567938
rect 366008 567854 366298 567882
rect 371634 567854 372016 567882
rect 376956 567868 376984 570687
rect 382094 570480 382150 570489
rect 382094 570415 382150 570424
rect 382108 567868 382136 570415
rect 392780 567868 392808 570959
rect 413926 570344 413982 570353
rect 408592 570308 408644 570314
rect 413926 570279 413982 570288
rect 408592 570250 408644 570256
rect 403254 570208 403310 570217
rect 403254 570143 403310 570152
rect 398104 568132 398156 568138
rect 398104 568074 398156 568080
rect 398116 567868 398144 568074
rect 403268 567868 403296 570143
rect 408604 567868 408632 570250
rect 413940 567868 413968 570279
rect 418724 567882 418752 576826
rect 424336 570654 424364 700334
rect 429856 699825 429884 703520
rect 439596 700868 439648 700874
rect 439596 700810 439648 700816
rect 439504 700732 439556 700738
rect 439504 700674 439556 700680
rect 429842 699816 429898 699825
rect 429842 699751 429898 699760
rect 439516 570790 439544 700674
rect 439504 570784 439556 570790
rect 439504 570726 439556 570732
rect 439608 570722 439636 700810
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 699718 494836 703520
rect 543476 700398 543504 703520
rect 559668 700534 559696 703520
rect 570328 700596 570380 700602
rect 570328 700538 570380 700544
rect 559656 700528 559708 700534
rect 559656 700470 559708 700476
rect 568856 700460 568908 700466
rect 568856 700402 568908 700408
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 568580 700392 568632 700398
rect 568580 700334 568632 700340
rect 494796 699712 494848 699718
rect 494796 699654 494848 699660
rect 495348 699712 495400 699718
rect 495348 699654 495400 699660
rect 495360 570790 495388 699654
rect 530216 570988 530268 570994
rect 530216 570930 530268 570936
rect 472072 570784 472124 570790
rect 472072 570726 472124 570732
rect 495348 570784 495400 570790
rect 495348 570726 495400 570732
rect 439596 570716 439648 570722
rect 439596 570658 439648 570664
rect 424324 570648 424376 570654
rect 424324 570590 424376 570596
rect 456248 570376 456300 570382
rect 456248 570318 456300 570324
rect 450912 570240 450964 570246
rect 450912 570182 450964 570188
rect 418724 567854 419106 567882
rect 424152 567866 424442 567882
rect 450924 567868 450952 570182
rect 456260 567868 456288 570318
rect 472084 567868 472112 570726
rect 519542 570616 519598 570625
rect 519542 570551 519598 570560
rect 477408 570172 477460 570178
rect 477408 570114 477460 570120
rect 477420 567868 477448 570114
rect 487896 570104 487948 570110
rect 487896 570046 487948 570052
rect 487908 567868 487936 570046
rect 509056 570036 509108 570042
rect 509056 569978 509108 569984
rect 509068 567868 509096 569978
rect 519556 567868 519584 570551
rect 524878 570072 524934 570081
rect 524878 570007 524934 570016
rect 524892 567868 524920 570007
rect 530228 567868 530256 570930
rect 535552 570784 535604 570790
rect 535552 570726 535604 570732
rect 535564 567868 535592 570726
rect 556712 570716 556764 570722
rect 556712 570658 556764 570664
rect 546038 570208 546094 570217
rect 546038 570143 546094 570152
rect 546052 567868 546080 570143
rect 556724 567868 556752 570658
rect 561864 570648 561916 570654
rect 561864 570590 561916 570596
rect 561876 567868 561904 570590
rect 424140 567860 424442 567866
rect 424192 567854 424442 567860
rect 424140 567802 424192 567808
rect 159732 567792 159784 567798
rect 202696 567792 202748 567798
rect 159784 567740 160034 567746
rect 159732 567734 160034 567740
rect 159744 567718 160034 567734
rect 202354 567740 202696 567746
rect 202354 567734 202748 567740
rect 202354 567718 202736 567734
rect 429488 567730 429778 567746
rect 429476 567724 429778 567730
rect 429528 567718 429778 567724
rect 429476 567666 429528 567672
rect 434812 567656 434864 567662
rect 445760 567656 445812 567662
rect 434864 567604 435114 567610
rect 434812 567598 435114 567604
rect 434824 567582 435114 567598
rect 445602 567604 445760 567610
rect 445602 567598 445812 567604
rect 445602 567582 445800 567598
rect 492968 567594 493258 567610
rect 492956 567588 493258 567594
rect 493008 567582 493258 567588
rect 492956 567530 493008 567536
rect 118056 567520 118108 567526
rect 112562 567458 112852 567474
rect 117714 567468 118056 567474
rect 117714 567462 118108 567468
rect 112562 567452 112864 567458
rect 112562 567446 112812 567452
rect 117714 567446 118096 567462
rect 112812 567394 112864 567400
rect 514116 567384 514168 567390
rect 86406 567352 86462 567361
rect 69952 567322 70242 567338
rect 69940 567316 70242 567322
rect 69992 567310 70242 567316
rect 86066 567310 86406 567338
rect 102046 567352 102102 567361
rect 91402 567322 91784 567338
rect 96554 567322 96752 567338
rect 91402 567316 91796 567322
rect 91402 567310 91744 567316
rect 86406 567287 86462 567296
rect 69940 567258 69992 567264
rect 96554 567316 96764 567322
rect 96554 567310 96712 567316
rect 91744 567258 91796 567264
rect 101890 567310 102046 567338
rect 128634 567352 128690 567361
rect 128386 567310 128634 567338
rect 102046 567287 102102 567296
rect 128634 567287 128690 567296
rect 133510 567352 133566 567361
rect 144550 567352 144606 567361
rect 133566 567310 133722 567338
rect 144210 567310 144550 567338
rect 133510 567287 133566 567296
rect 155222 567352 155278 567361
rect 154882 567310 155222 567338
rect 144550 567287 144606 567296
rect 170954 567352 171010 567361
rect 170706 567310 170954 567338
rect 155222 567287 155278 567296
rect 170954 567287 171010 567296
rect 212722 567352 212778 567361
rect 228546 567352 228602 567361
rect 212778 567310 213026 567338
rect 212722 567287 212778 567296
rect 244370 567352 244426 567361
rect 228602 567310 228850 567338
rect 228546 567287 228602 567296
rect 270866 567352 270922 567361
rect 244426 567310 244674 567338
rect 244370 567287 244426 567296
rect 281446 567352 281502 567361
rect 270922 567310 271170 567338
rect 270866 567287 270922 567296
rect 329010 567352 329066 567361
rect 281502 567310 281658 567338
rect 281446 567287 281502 567296
rect 339590 567352 339646 567361
rect 329066 567310 329314 567338
rect 329010 567287 329066 567296
rect 345294 567352 345350 567361
rect 339646 567310 339802 567338
rect 345138 567310 345294 567338
rect 339590 567287 339646 567296
rect 345294 567287 345350 567296
rect 387154 567352 387210 567361
rect 440054 567352 440110 567361
rect 387210 567310 387458 567338
rect 387154 567287 387210 567296
rect 461122 567352 461178 567361
rect 440110 567310 440266 567338
rect 440054 567287 440110 567296
rect 482282 567352 482338 567361
rect 461178 567310 461426 567338
rect 461122 567287 461178 567296
rect 482338 567310 482586 567338
rect 540426 567352 540482 567361
rect 514168 567332 514418 567338
rect 514116 567326 514418 567332
rect 514128 567310 514418 567326
rect 482282 567287 482338 567296
rect 551098 567352 551154 567361
rect 540482 567310 540730 567338
rect 540426 567287 540482 567296
rect 551154 567310 551402 567338
rect 567226 567310 567792 567338
rect 551098 567287 551154 567296
rect 96712 567258 96764 567264
rect 69848 310480 69900 310486
rect 69848 310422 69900 310428
rect 69848 247716 69900 247722
rect 69848 247658 69900 247664
rect 69756 3732 69808 3738
rect 69756 3674 69808 3680
rect 69860 3670 69888 247658
rect 70400 68740 70452 68746
rect 70400 68682 70452 68688
rect 132592 68740 132644 68746
rect 132592 68682 132644 68688
rect 153108 68740 153160 68746
rect 153108 68682 153160 68688
rect 70044 65074 70072 68068
rect 70032 65068 70084 65074
rect 70032 65010 70084 65016
rect 70412 16574 70440 68682
rect 72424 68604 72476 68610
rect 72424 68546 72476 68552
rect 128360 68604 128412 68610
rect 128360 68546 128412 68552
rect 71044 64252 71096 64258
rect 71044 64194 71096 64200
rect 70412 16546 70992 16574
rect 69848 3664 69900 3670
rect 69848 3606 69900 3612
rect 70308 3528 70360 3534
rect 70308 3470 70360 3476
rect 69572 3460 69624 3466
rect 69572 3402 69624 3408
rect 69112 2984 69164 2990
rect 69112 2926 69164 2932
rect 69124 480 69152 2926
rect 70320 480 70348 3470
rect 70964 3346 70992 16546
rect 71056 3534 71084 64194
rect 71688 7812 71740 7818
rect 71688 7754 71740 7760
rect 71044 3528 71096 3534
rect 71044 3470 71096 3476
rect 70964 3318 71544 3346
rect 71516 480 71544 3318
rect 71700 2990 71728 7754
rect 72436 3602 72464 68546
rect 84200 68536 84252 68542
rect 84200 68478 84252 68484
rect 126888 68536 126940 68542
rect 128372 68490 128400 68546
rect 126888 68478 126940 68484
rect 80152 68468 80204 68474
rect 80152 68410 80204 68416
rect 84108 68468 84160 68474
rect 84108 68410 84160 68416
rect 73160 68400 73212 68406
rect 73160 68342 73212 68348
rect 77208 68400 77260 68406
rect 77208 68342 77260 68348
rect 73068 68332 73120 68338
rect 73068 68274 73120 68280
rect 72424 3596 72476 3602
rect 72424 3538 72476 3544
rect 73080 3534 73108 68274
rect 73172 3534 73200 68342
rect 74632 67992 74684 67998
rect 74632 67934 74684 67940
rect 74644 16574 74672 67934
rect 75196 66094 75224 68068
rect 75184 66088 75236 66094
rect 75184 66030 75236 66036
rect 74644 16546 75040 16574
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73160 3528 73212 3534
rect 73160 3470 73212 3476
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 71688 2984 71740 2990
rect 71688 2926 71740 2932
rect 72620 480 72648 3470
rect 73816 480 73844 3470
rect 75012 480 75040 16546
rect 77220 3398 77248 68342
rect 79324 65408 79376 65414
rect 79324 65350 79376 65356
rect 77392 7608 77444 7614
rect 77392 7550 77444 7556
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 77208 3392 77260 3398
rect 77208 3334 77260 3340
rect 76208 480 76236 3334
rect 77404 480 77432 7550
rect 79336 3398 79364 65350
rect 79968 65000 80020 65006
rect 79968 64942 80020 64948
rect 79980 6914 80008 64942
rect 79704 6886 80008 6914
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 79324 3392 79376 3398
rect 79324 3334 79376 3340
rect 78600 480 78628 3334
rect 79704 480 79732 6886
rect 80164 3398 80192 68410
rect 80532 66094 80560 68068
rect 80520 66088 80572 66094
rect 80520 66030 80572 66036
rect 81348 66088 81400 66094
rect 81348 66030 81400 66036
rect 81360 5370 81388 66030
rect 81440 65068 81492 65074
rect 81440 65010 81492 65016
rect 81452 16574 81480 65010
rect 81452 16546 81664 16574
rect 81348 5364 81400 5370
rect 81348 5306 81400 5312
rect 80152 3392 80204 3398
rect 80152 3334 80204 3340
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 80900 480 80928 3334
rect 81636 490 81664 16546
rect 84120 3398 84148 68410
rect 84212 16574 84240 68478
rect 85868 65754 85896 68068
rect 90744 68054 91034 68082
rect 96370 68054 96568 68082
rect 101706 68054 102088 68082
rect 90744 66230 90772 68054
rect 91100 67040 91152 67046
rect 91100 66982 91152 66988
rect 90732 66224 90784 66230
rect 90732 66166 90784 66172
rect 91008 66224 91060 66230
rect 91008 66166 91060 66172
rect 85856 65748 85908 65754
rect 85856 65690 85908 65696
rect 84212 16546 84516 16574
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 81912 598 82124 626
rect 81912 490 81940 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 462 81940 490
rect 82096 480 82124 598
rect 83292 480 83320 3334
rect 84488 480 84516 16546
rect 86868 5228 86920 5234
rect 86868 5170 86920 5176
rect 85672 3460 85724 3466
rect 85672 3402 85724 3408
rect 85684 480 85712 3402
rect 86880 480 86908 5170
rect 91020 3534 91048 66166
rect 91112 16574 91140 66982
rect 95148 65748 95200 65754
rect 95148 65690 95200 65696
rect 91112 16546 91600 16574
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 87972 3460 88024 3466
rect 87972 3402 88024 3408
rect 87984 480 88012 3402
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 16546
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 93952 3528 94004 3534
rect 92754 3496 92810 3505
rect 93952 3470 94004 3476
rect 92754 3431 92810 3440
rect 92768 480 92796 3431
rect 93964 480 93992 3470
rect 95068 1850 95096 3538
rect 95160 3534 95188 65690
rect 96540 5302 96568 68054
rect 100668 65068 100720 65074
rect 100668 65010 100720 65016
rect 96252 5296 96304 5302
rect 96252 5238 96304 5244
rect 96528 5296 96580 5302
rect 96528 5238 96580 5244
rect 95148 3528 95200 3534
rect 95148 3470 95200 3476
rect 95068 1822 95188 1850
rect 95160 480 95188 1822
rect 96264 480 96292 5238
rect 98644 4072 98696 4078
rect 98644 4014 98696 4020
rect 97446 3496 97502 3505
rect 97446 3431 97502 3440
rect 97460 480 97488 3431
rect 98656 480 98684 4014
rect 100680 3534 100708 65010
rect 102060 64874 102088 68054
rect 107028 66026 107056 68068
rect 111708 67040 111760 67046
rect 111708 66982 111760 66988
rect 107016 66020 107068 66026
rect 107016 65962 107068 65968
rect 104808 65000 104860 65006
rect 104808 64942 104860 64948
rect 102060 64846 102272 64874
rect 102244 16574 102272 64846
rect 102244 16546 103376 16574
rect 101036 6180 101088 6186
rect 101036 6122 101088 6128
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 99852 480 99880 3470
rect 101048 480 101076 6122
rect 102232 3392 102284 3398
rect 102232 3334 102284 3340
rect 102244 480 102272 3334
rect 103348 480 103376 16546
rect 104820 6914 104848 64942
rect 111720 6914 111748 66982
rect 112180 65006 112208 68068
rect 117332 68054 117530 68082
rect 115848 67108 115900 67114
rect 115848 67050 115900 67056
rect 112168 65000 112220 65006
rect 112168 64942 112220 64948
rect 113088 65000 113140 65006
rect 113088 64942 113140 64948
rect 113100 6914 113128 64942
rect 104544 6886 104848 6914
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 104544 480 104572 6886
rect 109314 5264 109370 5273
rect 109314 5199 109370 5208
rect 108118 4992 108174 5001
rect 108118 4927 108174 4936
rect 106922 3632 106978 3641
rect 106922 3567 106978 3576
rect 105726 3360 105782 3369
rect 105726 3295 105782 3304
rect 105740 480 105768 3295
rect 106936 480 106964 3567
rect 108132 480 108160 4927
rect 109328 480 109356 5199
rect 110510 3496 110566 3505
rect 110510 3431 110566 3440
rect 110524 480 110552 3431
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114008 4072 114060 4078
rect 114008 4014 114060 4020
rect 114020 480 114048 4014
rect 115860 3602 115888 67050
rect 117332 64326 117360 68054
rect 119988 67176 120040 67182
rect 119988 67118 120040 67124
rect 117320 64320 117372 64326
rect 117320 64262 117372 64268
rect 120000 6914 120028 67118
rect 122748 64184 122800 64190
rect 122748 64126 122800 64132
rect 119908 6886 120028 6914
rect 118790 4856 118846 4865
rect 118790 4791 118846 4800
rect 117594 3632 117650 3641
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 116400 3596 116452 3602
rect 117594 3567 117650 3576
rect 116400 3538 116452 3544
rect 115216 480 115244 3538
rect 116412 480 116440 3538
rect 117608 480 117636 3567
rect 118804 480 118832 4791
rect 119908 480 119936 6886
rect 121092 3732 121144 3738
rect 121092 3674 121144 3680
rect 121104 480 121132 3674
rect 122760 3398 122788 64126
rect 123484 3664 123536 3670
rect 123484 3606 123536 3612
rect 124680 3664 124732 3670
rect 124680 3606 124732 3612
rect 122288 3392 122340 3398
rect 122288 3334 122340 3340
rect 122748 3392 122800 3398
rect 122748 3334 122800 3340
rect 122300 480 122328 3334
rect 123496 480 123524 3606
rect 124692 480 124720 3606
rect 126900 3398 126928 68478
rect 128280 68462 128400 68490
rect 128188 67250 128216 68068
rect 128176 67244 128228 67250
rect 128176 67186 128228 67192
rect 128176 5364 128228 5370
rect 128176 5306 128228 5312
rect 125876 3392 125928 3398
rect 125876 3334 125928 3340
rect 126888 3392 126940 3398
rect 126888 3334 126940 3340
rect 126980 3392 127032 3398
rect 126980 3334 127032 3340
rect 125888 480 125916 3334
rect 126992 480 127020 3334
rect 128188 480 128216 5306
rect 128280 3398 128308 68462
rect 130384 66020 130436 66026
rect 130384 65962 130436 65968
rect 128360 64388 128412 64394
rect 128360 64330 128412 64336
rect 128372 16574 128400 64330
rect 128372 16546 128952 16574
rect 128268 3392 128320 3398
rect 128268 3334 128320 3340
rect 128924 490 128952 16546
rect 130396 4894 130424 65962
rect 132604 16574 132632 68682
rect 140780 68672 140832 68678
rect 140780 68614 140832 68620
rect 133340 65346 133368 68068
rect 138032 68054 138690 68082
rect 133328 65340 133380 65346
rect 133328 65282 133380 65288
rect 138032 64394 138060 68054
rect 138020 64388 138072 64394
rect 138020 64330 138072 64336
rect 140792 16574 140820 68614
rect 144012 65346 144040 68068
rect 149072 68054 149362 68082
rect 144000 65340 144052 65346
rect 144000 65282 144052 65288
rect 144828 65340 144880 65346
rect 144828 65282 144880 65288
rect 144736 18624 144788 18630
rect 144736 18566 144788 18572
rect 132604 16546 133000 16574
rect 140792 16546 141280 16574
rect 131764 7676 131816 7682
rect 131764 7618 131816 7624
rect 130384 4888 130436 4894
rect 130384 4830 130436 4836
rect 130566 3768 130622 3777
rect 130566 3703 130622 3712
rect 129200 598 129412 626
rect 129200 490 129228 598
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 462 129228 490
rect 129384 480 129412 598
rect 130580 480 130608 3703
rect 131776 480 131804 7618
rect 132972 480 133000 16546
rect 134156 6860 134208 6866
rect 134156 6802 134208 6808
rect 134168 480 134196 6802
rect 138848 6520 138900 6526
rect 138848 6462 138900 6468
rect 135258 5128 135314 5137
rect 135258 5063 135314 5072
rect 135272 480 135300 5063
rect 137652 4956 137704 4962
rect 137652 4898 137704 4904
rect 136456 4888 136508 4894
rect 136456 4830 136508 4836
rect 136468 480 136496 4830
rect 137664 480 137692 4898
rect 138860 480 138888 6462
rect 140042 3768 140098 3777
rect 140042 3703 140098 3712
rect 140056 480 140084 3703
rect 141252 480 141280 16546
rect 142436 6588 142488 6594
rect 142436 6530 142488 6536
rect 142448 480 142476 6530
rect 143540 4956 143592 4962
rect 143540 4898 143592 4904
rect 143552 480 143580 4898
rect 144748 480 144776 18566
rect 144840 6322 144868 65282
rect 149072 20670 149100 68054
rect 150348 67652 150400 67658
rect 150348 67594 150400 67600
rect 149060 20664 149112 20670
rect 149060 20606 149112 20612
rect 148324 6452 148376 6458
rect 148324 6394 148376 6400
rect 144828 6316 144880 6322
rect 144828 6258 144880 6264
rect 147128 6248 147180 6254
rect 147128 6190 147180 6196
rect 145930 3768 145986 3777
rect 145930 3703 145986 3712
rect 145944 480 145972 3703
rect 147140 480 147168 6190
rect 148336 480 148364 6394
rect 150360 3398 150388 67594
rect 150622 6760 150678 6769
rect 150622 6695 150678 6704
rect 149520 3392 149572 3398
rect 149520 3334 149572 3340
rect 150348 3392 150400 3398
rect 150348 3334 150400 3340
rect 149532 480 149560 3334
rect 150636 480 150664 6695
rect 153014 3768 153070 3777
rect 153014 3703 153070 3712
rect 151820 3392 151872 3398
rect 151820 3334 151872 3340
rect 151832 480 151860 3334
rect 153028 480 153056 3703
rect 153120 3398 153148 68682
rect 190552 68264 190604 68270
rect 190552 68206 190604 68212
rect 197360 68264 197412 68270
rect 197360 68206 197412 68212
rect 200028 68264 200080 68270
rect 200028 68206 200080 68212
rect 206928 68264 206980 68270
rect 206928 68206 206980 68212
rect 154304 67652 154356 67658
rect 154304 67594 154356 67600
rect 154316 6914 154344 67594
rect 154500 65074 154528 68068
rect 159284 68054 159850 68082
rect 157340 67720 157392 67726
rect 157340 67662 157392 67668
rect 154488 65068 154540 65074
rect 154488 65010 154540 65016
rect 157352 16574 157380 67662
rect 159284 65890 159312 68054
rect 161480 67788 161532 67794
rect 161480 67730 161532 67736
rect 159272 65884 159324 65890
rect 159272 65826 159324 65832
rect 159364 65884 159416 65890
rect 159364 65826 159416 65832
rect 158720 62824 158772 62830
rect 158720 62766 158772 62772
rect 158732 16574 158760 62766
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 154224 6886 154344 6914
rect 153108 3392 153160 3398
rect 153108 3334 153160 3340
rect 154224 480 154252 6886
rect 155408 6384 155460 6390
rect 155408 6326 155460 6332
rect 155420 480 155448 6326
rect 156602 3768 156658 3777
rect 156602 3703 156658 3712
rect 156616 480 156644 3703
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 159376 6526 159404 65826
rect 160744 65340 160796 65346
rect 160744 65282 160796 65288
rect 160756 6594 160784 65282
rect 161492 16574 161520 67730
rect 165172 65890 165200 68068
rect 167000 67856 167052 67862
rect 167000 67798 167052 67804
rect 165160 65884 165212 65890
rect 165160 65826 165212 65832
rect 162860 64388 162912 64394
rect 162860 64330 162912 64336
rect 162872 16574 162900 64330
rect 167012 16574 167040 67798
rect 175660 66842 175688 68068
rect 178040 67856 178092 67862
rect 178040 67798 178092 67804
rect 175648 66836 175700 66842
rect 175648 66778 175700 66784
rect 168380 66632 168432 66638
rect 168380 66574 168432 66580
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 167012 16546 167224 16574
rect 160744 6588 160796 6594
rect 160744 6530 160796 6536
rect 159364 6520 159416 6526
rect 159364 6462 159416 6468
rect 161294 5944 161350 5953
rect 161294 5879 161350 5888
rect 160098 3768 160154 3777
rect 160098 3703 160154 3712
rect 160112 480 160140 3703
rect 161308 480 161336 5879
rect 162044 490 162072 16546
rect 162320 598 162532 626
rect 162320 490 162348 598
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 462 162348 490
rect 162504 480 162532 598
rect 163700 480 163728 16546
rect 166078 5536 166134 5545
rect 166078 5471 166134 5480
rect 164882 3768 164938 3777
rect 164882 3703 164938 3712
rect 164896 480 164924 3703
rect 166092 480 166120 5471
rect 167196 480 167224 16546
rect 168392 11762 168420 66574
rect 175280 57248 175332 57254
rect 175280 57190 175332 57196
rect 175292 16574 175320 57190
rect 178052 16574 178080 67798
rect 180996 67289 181024 68068
rect 182180 67856 182232 67862
rect 182180 67798 182232 67804
rect 186044 67856 186096 67862
rect 186044 67798 186096 67804
rect 190368 67856 190420 67862
rect 190368 67798 190420 67804
rect 180982 67280 181038 67289
rect 180982 67215 181038 67224
rect 181444 65068 181496 65074
rect 181444 65010 181496 65016
rect 175292 16546 175504 16574
rect 178052 16546 178632 16574
rect 168380 11756 168432 11762
rect 168380 11698 168432 11704
rect 169576 11756 169628 11762
rect 169576 11698 169628 11704
rect 168378 5128 168434 5137
rect 168378 5063 168434 5072
rect 168392 480 168420 5063
rect 169588 480 169616 11698
rect 174268 6588 174320 6594
rect 174268 6530 174320 6536
rect 173164 6316 173216 6322
rect 173164 6258 173216 6264
rect 171968 5024 172020 5030
rect 170770 4992 170826 5001
rect 171968 4966 172020 4972
rect 170770 4927 170826 4936
rect 170784 480 170812 4927
rect 171980 480 172008 4966
rect 173176 480 173204 6258
rect 174280 480 174308 6530
rect 175476 480 175504 16546
rect 176660 6792 176712 6798
rect 176660 6734 176712 6740
rect 176672 480 176700 6734
rect 177856 5024 177908 5030
rect 177856 4966 177908 4972
rect 177868 480 177896 4966
rect 178604 490 178632 16546
rect 180246 6216 180302 6225
rect 181456 6186 181484 65010
rect 181536 6656 181588 6662
rect 181536 6598 181588 6604
rect 180246 6151 180302 6160
rect 181444 6180 181496 6186
rect 178880 598 179092 626
rect 178880 490 178908 598
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 462 178908 490
rect 179064 480 179092 598
rect 180260 480 180288 6151
rect 181444 6122 181496 6128
rect 181548 3346 181576 6598
rect 181456 3318 181576 3346
rect 181456 480 181484 3318
rect 182192 490 182220 67798
rect 184204 65884 184256 65890
rect 184204 65826 184256 65832
rect 183742 6080 183798 6089
rect 183742 6015 183798 6024
rect 182376 598 182588 626
rect 182376 490 182404 598
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 462 182404 490
rect 182560 480 182588 598
rect 183756 480 183784 6015
rect 184216 3670 184244 65826
rect 184204 3664 184256 3670
rect 184204 3606 184256 3612
rect 186056 3398 186084 67798
rect 187700 66700 187752 66706
rect 187700 66642 187752 66648
rect 187712 16574 187740 66642
rect 187712 16546 188568 16574
rect 186136 6520 186188 6526
rect 186136 6462 186188 6468
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 186044 3392 186096 3398
rect 186044 3334 186096 3340
rect 184952 480 184980 3334
rect 186148 480 186176 6462
rect 187332 6180 187384 6186
rect 187332 6122 187384 6128
rect 187344 480 187372 6122
rect 188540 480 188568 16546
rect 190380 3398 190408 67798
rect 190564 16574 190592 68206
rect 191484 65142 191512 68068
rect 191472 65136 191524 65142
rect 191472 65078 191524 65084
rect 196820 65006 196848 68068
rect 196808 65000 196860 65006
rect 196808 64942 196860 64948
rect 197268 64388 197320 64394
rect 197268 64330 197320 64336
rect 194508 62824 194560 62830
rect 194508 62766 194560 62772
rect 190564 16546 190868 16574
rect 189724 3392 189776 3398
rect 189724 3334 189776 3340
rect 190368 3392 190420 3398
rect 190368 3334 190420 3340
rect 189736 480 189764 3334
rect 190840 480 190868 16546
rect 194520 6914 194548 62766
rect 194428 6886 194548 6914
rect 192024 6724 192076 6730
rect 192024 6666 192076 6672
rect 192036 480 192064 6666
rect 193220 5296 193272 5302
rect 193220 5238 193272 5244
rect 193232 480 193260 5238
rect 194428 480 194456 6886
rect 195610 6352 195666 6361
rect 195610 6287 195666 6296
rect 195624 480 195652 6287
rect 197280 3398 197308 64330
rect 197372 16574 197400 68206
rect 197372 16546 197952 16574
rect 196808 3392 196860 3398
rect 196808 3334 196860 3340
rect 197268 3392 197320 3398
rect 197268 3334 197320 3340
rect 196820 480 196848 3334
rect 197924 480 197952 16546
rect 200040 3398 200068 68206
rect 202170 68054 202828 68082
rect 202696 46232 202748 46238
rect 202696 46174 202748 46180
rect 200302 6624 200358 6633
rect 200302 6559 200358 6568
rect 199108 3392 199160 3398
rect 199108 3334 199160 3340
rect 200028 3392 200080 3398
rect 200028 3334 200080 3340
rect 199120 480 199148 3334
rect 200316 480 200344 6559
rect 201498 5400 201554 5409
rect 201498 5335 201554 5344
rect 201512 480 201540 5335
rect 202708 480 202736 46174
rect 202800 20670 202828 68054
rect 202788 20664 202840 20670
rect 202788 20606 202840 20612
rect 203890 5264 203946 5273
rect 203890 5199 203946 5208
rect 203904 480 203932 5199
rect 205086 3632 205142 3641
rect 205086 3567 205142 3576
rect 205100 480 205128 3567
rect 206940 3398 206968 68206
rect 211160 68196 211212 68202
rect 211160 68138 211212 68144
rect 219348 68196 219400 68202
rect 219348 68138 219400 68144
rect 207032 68054 207506 68082
rect 207032 5030 207060 68054
rect 209780 67924 209832 67930
rect 209780 67866 209832 67872
rect 208400 66768 208452 66774
rect 208400 66710 208452 66716
rect 208412 16574 208440 66710
rect 208412 16546 208624 16574
rect 207020 5024 207072 5030
rect 207020 4966 207072 4972
rect 207388 5024 207440 5030
rect 207388 4966 207440 4972
rect 206192 3392 206244 3398
rect 206192 3334 206244 3340
rect 206928 3392 206980 3398
rect 206928 3334 206980 3340
rect 206204 480 206232 3334
rect 207400 480 207428 4966
rect 208596 480 208624 16546
rect 209792 480 209820 67866
rect 211172 16574 211200 68138
rect 217980 65278 218008 68068
rect 217968 65272 218020 65278
rect 217968 65214 218020 65220
rect 211172 16546 211752 16574
rect 210974 3632 211030 3641
rect 210974 3567 211030 3576
rect 210988 480 211016 3567
rect 211724 490 211752 16546
rect 216864 7744 216916 7750
rect 216864 7686 216916 7692
rect 214472 5092 214524 5098
rect 214472 5034 214524 5040
rect 213368 3664 213420 3670
rect 213368 3606 213420 3612
rect 212000 598 212212 626
rect 212000 490 212028 598
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 462 212028 490
rect 212184 480 212212 598
rect 213380 480 213408 3606
rect 214484 480 214512 5034
rect 215668 3732 215720 3738
rect 215668 3674 215720 3680
rect 215680 480 215708 3674
rect 216876 480 216904 7686
rect 219256 6316 219308 6322
rect 219256 6258 219308 6264
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218072 480 218100 3334
rect 219268 480 219296 6258
rect 219360 3398 219388 68138
rect 222200 68128 222252 68134
rect 222200 68070 222252 68076
rect 226248 68128 226300 68134
rect 226248 68070 226300 68076
rect 220820 67992 220872 67998
rect 220820 67934 220872 67940
rect 220832 16574 220860 67934
rect 222212 16574 222240 68070
rect 223316 67561 223344 68068
rect 223302 67552 223358 67561
rect 223302 67487 223358 67496
rect 224868 65136 224920 65142
rect 224868 65078 224920 65084
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 220450 3632 220506 3641
rect 220450 3567 220506 3576
rect 219348 3392 219400 3398
rect 219348 3334 219400 3340
rect 220464 480 220492 3567
rect 221108 490 221136 16546
rect 221384 598 221596 626
rect 221384 490 221412 598
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 462 221412 490
rect 221568 480 221596 598
rect 222764 480 222792 16546
rect 224880 3398 224908 65078
rect 226260 3398 226288 68070
rect 227812 68060 227864 68066
rect 227812 68002 227864 68008
rect 227824 16574 227852 68002
rect 228652 65210 228680 68068
rect 230388 68060 230440 68066
rect 230388 68002 230440 68008
rect 238772 68054 239154 68082
rect 244292 68054 244490 68082
rect 228640 65204 228692 65210
rect 228640 65146 228692 65152
rect 227824 16546 228312 16574
rect 226338 6896 226394 6905
rect 226338 6831 226394 6840
rect 223948 3392 224000 3398
rect 223948 3334 224000 3340
rect 224868 3392 224920 3398
rect 224868 3334 224920 3340
rect 225144 3392 225196 3398
rect 225144 3334 225196 3340
rect 226248 3392 226300 3398
rect 226248 3334 226300 3340
rect 223960 480 223988 3334
rect 225156 480 225184 3334
rect 226352 480 226380 6831
rect 227534 3632 227590 3641
rect 227534 3567 227590 3576
rect 227548 480 227576 3567
rect 228284 490 228312 16546
rect 230400 3398 230428 68002
rect 235816 65272 235868 65278
rect 235816 65214 235868 65220
rect 230480 64320 230532 64326
rect 230480 64262 230532 64268
rect 230492 16574 230520 64262
rect 230492 16546 231072 16574
rect 229836 3392 229888 3398
rect 229836 3334 229888 3340
rect 230388 3392 230440 3398
rect 230388 3334 230440 3340
rect 228560 598 228772 626
rect 228560 490 228588 598
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 462 228588 490
rect 228744 480 228772 598
rect 229848 480 229876 3334
rect 231044 480 231072 16546
rect 233422 6488 233478 6497
rect 233422 6423 233478 6432
rect 232228 5296 232280 5302
rect 232228 5238 232280 5244
rect 232240 480 232268 5238
rect 233436 480 233464 6423
rect 235828 3398 235856 65214
rect 238772 64394 238800 68054
rect 238760 64388 238812 64394
rect 238760 64330 238812 64336
rect 244292 6866 244320 68054
rect 249812 18630 249840 68068
rect 254964 66842 254992 68068
rect 254952 66836 255004 66842
rect 254952 66778 255004 66784
rect 260300 66774 260328 68068
rect 270512 68054 270986 68082
rect 260288 66768 260340 66774
rect 260288 66710 260340 66716
rect 249800 18624 249852 18630
rect 249800 18566 249852 18572
rect 244280 6860 244332 6866
rect 244280 6802 244332 6808
rect 237010 6488 237066 6497
rect 237010 6423 237066 6432
rect 235908 5092 235960 5098
rect 235908 5034 235960 5040
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 234632 480 234660 3334
rect 235920 2530 235948 5034
rect 235828 2502 235948 2530
rect 235828 480 235856 2502
rect 237024 480 237052 6423
rect 270512 5166 270540 68054
rect 276124 65278 276152 68068
rect 276112 65272 276164 65278
rect 276112 65214 276164 65220
rect 276664 65272 276716 65278
rect 276664 65214 276716 65220
rect 270500 5160 270552 5166
rect 238114 5128 238170 5137
rect 270500 5102 270552 5108
rect 238114 5063 238170 5072
rect 238128 480 238156 5063
rect 276676 4010 276704 65214
rect 280804 65204 280856 65210
rect 280804 65146 280856 65152
rect 276664 4004 276716 4010
rect 276664 3946 276716 3952
rect 280816 3874 280844 65146
rect 281460 65074 281488 68068
rect 285692 68054 286810 68082
rect 281448 65068 281500 65074
rect 281448 65010 281500 65016
rect 285692 5234 285720 68054
rect 292132 65074 292160 68068
rect 296732 68054 297298 68082
rect 286324 65068 286376 65074
rect 286324 65010 286376 65016
rect 292120 65068 292172 65074
rect 292120 65010 292172 65016
rect 285680 5228 285732 5234
rect 285680 5170 285732 5176
rect 286336 4078 286364 65010
rect 291844 65000 291896 65006
rect 291844 64942 291896 64948
rect 286324 4072 286376 4078
rect 286324 4014 286376 4020
rect 291856 3942 291884 64942
rect 296732 64258 296760 68054
rect 307956 67425 307984 68068
rect 311912 68054 313122 68082
rect 307942 67416 307998 67425
rect 307942 67351 307998 67360
rect 297364 65068 297416 65074
rect 297364 65010 297416 65016
rect 296720 64252 296772 64258
rect 296720 64194 296772 64200
rect 291844 3936 291896 3942
rect 291844 3878 291896 3884
rect 280804 3868 280856 3874
rect 280804 3810 280856 3816
rect 297376 3806 297404 65010
rect 311912 7818 311940 68054
rect 318444 65006 318472 68068
rect 323780 65482 323808 68068
rect 329116 66706 329144 68068
rect 333992 68054 334282 68082
rect 329104 66700 329156 66706
rect 329104 66642 329156 66648
rect 323768 65476 323820 65482
rect 323768 65418 323820 65424
rect 318432 65000 318484 65006
rect 318432 64942 318484 64948
rect 311900 7812 311952 7818
rect 311900 7754 311952 7760
rect 333992 6798 334020 68054
rect 339604 64874 339632 68068
rect 344940 65414 344968 68068
rect 349172 68054 350290 68082
rect 345664 65476 345716 65482
rect 345664 65418 345716 65424
rect 344928 65408 344980 65414
rect 344928 65350 344980 65356
rect 339512 64846 339632 64874
rect 333980 6792 334032 6798
rect 333980 6734 334032 6740
rect 339512 6662 339540 64846
rect 339500 6656 339552 6662
rect 339500 6598 339552 6604
rect 345676 6594 345704 65418
rect 349172 6730 349200 68054
rect 355428 65482 355456 68068
rect 360764 66162 360792 68068
rect 366100 67250 366128 68068
rect 366088 67244 366140 67250
rect 366088 67186 366140 67192
rect 360752 66156 360804 66162
rect 360752 66098 360804 66104
rect 355416 65476 355468 65482
rect 355416 65418 355468 65424
rect 371436 65074 371464 68068
rect 376588 66570 376616 68068
rect 376576 66564 376628 66570
rect 376576 66506 376628 66512
rect 381924 66230 381952 68068
rect 387260 67318 387288 68068
rect 387248 67312 387300 67318
rect 387248 67254 387300 67260
rect 381912 66224 381964 66230
rect 381912 66166 381964 66172
rect 371884 66156 371936 66162
rect 371884 66098 371936 66104
rect 371424 65068 371476 65074
rect 371424 65010 371476 65016
rect 349160 6724 349212 6730
rect 349160 6666 349212 6672
rect 345664 6588 345716 6594
rect 345664 6530 345716 6536
rect 371896 6526 371924 66098
rect 392596 65210 392624 68068
rect 397748 65958 397776 68068
rect 403084 66230 403112 68068
rect 403072 66224 403124 66230
rect 403072 66166 403124 66172
rect 397736 65952 397788 65958
rect 397736 65894 397788 65900
rect 392584 65204 392636 65210
rect 392584 65146 392636 65152
rect 408420 65142 408448 68068
rect 412652 68054 413586 68082
rect 408408 65136 408460 65142
rect 408408 65078 408460 65084
rect 371884 6520 371936 6526
rect 371884 6462 371936 6468
rect 412652 5302 412680 68054
rect 418908 67386 418936 68068
rect 418896 67380 418948 67386
rect 418896 67322 418948 67328
rect 424244 65346 424272 68068
rect 429212 68054 429594 68082
rect 424232 65340 424284 65346
rect 424232 65282 424284 65288
rect 429212 7682 429240 68054
rect 429200 7676 429252 7682
rect 429200 7618 429252 7624
rect 434732 6458 434760 68068
rect 440068 66094 440096 68068
rect 450740 66094 450768 68068
rect 455432 68054 455906 68082
rect 440056 66088 440108 66094
rect 440056 66030 440108 66036
rect 450728 66088 450780 66094
rect 450728 66030 450780 66036
rect 434720 6452 434772 6458
rect 434720 6394 434772 6400
rect 412640 5296 412692 5302
rect 412640 5238 412692 5244
rect 455432 5030 455460 68054
rect 461228 65822 461256 68068
rect 461216 65816 461268 65822
rect 461216 65758 461268 65764
rect 466564 64874 466592 68068
rect 466472 64846 466592 64874
rect 470612 68054 471914 68082
rect 466472 6390 466500 64846
rect 470612 7750 470640 68054
rect 477052 67454 477080 68068
rect 481652 68054 482402 68082
rect 477040 67448 477092 67454
rect 477040 67390 477092 67396
rect 470600 7744 470652 7750
rect 470600 7686 470652 7692
rect 466460 6384 466512 6390
rect 466460 6326 466512 6332
rect 481652 5098 481680 68054
rect 487724 65618 487752 68068
rect 498212 65686 498240 68068
rect 503548 67522 503576 68068
rect 503536 67516 503588 67522
rect 503536 67458 503588 67464
rect 508884 66026 508912 68068
rect 518912 68054 519386 68082
rect 508872 66020 508924 66026
rect 508872 65962 508924 65968
rect 498200 65680 498252 65686
rect 498200 65622 498252 65628
rect 487712 65612 487764 65618
rect 487712 65554 487764 65560
rect 518912 6254 518940 68054
rect 524708 65278 524736 68068
rect 535196 66162 535224 68068
rect 535184 66156 535236 66162
rect 535184 66098 535236 66104
rect 540532 65754 540560 68068
rect 545868 67590 545896 68068
rect 550652 68054 551218 68082
rect 545856 67584 545908 67590
rect 545856 67526 545908 67532
rect 540520 65748 540572 65754
rect 540520 65690 540572 65696
rect 524696 65272 524748 65278
rect 524696 65214 524748 65220
rect 518900 6248 518952 6254
rect 518900 6190 518952 6196
rect 481640 5092 481692 5098
rect 481640 5034 481692 5040
rect 455420 5024 455472 5030
rect 455420 4966 455472 4972
rect 550652 4962 550680 68054
rect 567028 65550 567056 68068
rect 567016 65544 567068 65550
rect 567016 65486 567068 65492
rect 567764 46238 567792 567310
rect 568592 565962 568620 700334
rect 568764 566024 568816 566030
rect 568764 565966 568816 565972
rect 568580 565956 568632 565962
rect 568580 565898 568632 565904
rect 568776 540974 568804 565966
rect 568500 540946 568804 540974
rect 568500 525794 568528 540946
rect 568868 540274 568896 700402
rect 570052 700324 570104 700330
rect 570052 700266 570104 700272
rect 569960 683188 570012 683194
rect 569960 683130 570012 683136
rect 569316 570308 569368 570314
rect 569316 570250 569368 570256
rect 568948 548140 569000 548146
rect 568948 548082 569000 548088
rect 568960 540394 568988 548082
rect 568948 540388 569000 540394
rect 568948 540330 569000 540336
rect 568868 540246 569080 540274
rect 568408 525766 568528 525794
rect 568408 497944 568436 525766
rect 568948 525360 569000 525366
rect 568500 525308 568948 525314
rect 568500 525302 569000 525308
rect 568500 525286 568988 525302
rect 568500 516202 568528 525286
rect 569052 516202 569080 540246
rect 568500 516174 568620 516202
rect 568592 516134 568620 516174
rect 568868 516174 569080 516202
rect 568592 516106 568804 516134
rect 568776 503146 568804 516106
rect 568868 507854 568896 516174
rect 568868 507826 568988 507854
rect 568776 503118 568896 503146
rect 568868 502334 568896 503118
rect 568960 503062 568988 507826
rect 568948 503056 569000 503062
rect 568948 502998 569000 503004
rect 568868 502306 568988 502334
rect 568960 498098 568988 502306
rect 569040 499792 569092 499798
rect 569040 499734 569092 499740
rect 568948 498092 569000 498098
rect 568948 498034 569000 498040
rect 568948 497956 569000 497962
rect 568408 497916 568948 497944
rect 568948 497898 569000 497904
rect 568948 497820 569000 497826
rect 568948 497762 569000 497768
rect 568960 497570 568988 497762
rect 568592 497542 568988 497570
rect 567844 69828 567896 69834
rect 567844 69770 567896 69776
rect 567752 46232 567804 46238
rect 567752 46174 567804 46180
rect 550640 4956 550692 4962
rect 550640 4898 550692 4904
rect 297364 3800 297416 3806
rect 297364 3742 297416 3748
rect 567856 3602 567884 69770
rect 568592 7614 568620 497542
rect 568948 495372 569000 495378
rect 568948 495314 569000 495320
rect 568960 492674 568988 495314
rect 568684 492646 568988 492674
rect 568684 491294 568712 492646
rect 568684 491266 568988 491294
rect 568960 486470 568988 491266
rect 568948 486464 569000 486470
rect 568948 486406 569000 486412
rect 569052 486146 569080 499734
rect 568684 486118 569080 486146
rect 568684 68474 568712 486118
rect 568948 485104 569000 485110
rect 568948 485046 569000 485052
rect 568960 481634 568988 485046
rect 568868 481606 568988 481634
rect 568868 460934 568896 481606
rect 568868 460906 569080 460934
rect 568948 445800 569000 445806
rect 568948 445742 569000 445748
rect 568960 444258 568988 445742
rect 568776 444230 568988 444258
rect 568672 68468 568724 68474
rect 568672 68410 568724 68416
rect 568776 67114 568804 444230
rect 569052 441674 569080 460906
rect 568868 441646 569080 441674
rect 568868 441614 568896 441646
rect 568868 441586 568988 441614
rect 568960 431594 568988 441586
rect 568948 431588 569000 431594
rect 568948 431530 569000 431536
rect 569224 390584 569276 390590
rect 569224 390526 569276 390532
rect 568948 321632 569000 321638
rect 568948 321574 569000 321580
rect 568960 316034 568988 321574
rect 568868 316006 568988 316034
rect 568764 67108 568816 67114
rect 568764 67050 568816 67056
rect 568580 7608 568632 7614
rect 568580 7550 568632 7556
rect 568868 3738 568896 316006
rect 569040 266416 569092 266422
rect 569040 266358 569092 266364
rect 568948 219768 569000 219774
rect 568948 219710 569000 219716
rect 568960 4826 568988 219710
rect 569052 69358 569080 266358
rect 569132 258528 569184 258534
rect 569132 258470 569184 258476
rect 569040 69352 569092 69358
rect 569040 69294 569092 69300
rect 569144 68066 569172 258470
rect 569132 68060 569184 68066
rect 569132 68002 569184 68008
rect 568948 4820 569000 4826
rect 568948 4762 569000 4768
rect 568856 3732 568908 3738
rect 568856 3674 568908 3680
rect 567844 3596 567896 3602
rect 567844 3538 567896 3544
rect 569236 3466 569264 390526
rect 569328 365702 569356 570250
rect 569408 565956 569460 565962
rect 569408 565898 569460 565904
rect 569420 564369 569448 565898
rect 569406 564360 569462 564369
rect 569406 564295 569462 564304
rect 569406 548176 569462 548185
rect 569406 548111 569408 548120
rect 569460 548111 569462 548120
rect 569408 548082 569460 548088
rect 569406 500848 569462 500857
rect 569406 500783 569462 500792
rect 569420 499798 569448 500783
rect 569408 499792 569460 499798
rect 569408 499734 569460 499740
rect 569408 497956 569460 497962
rect 569408 497898 569460 497904
rect 569420 494057 569448 497898
rect 569406 494048 569462 494057
rect 569406 493983 569462 493992
rect 569406 446176 569462 446185
rect 569406 446111 569462 446120
rect 569420 445806 569448 446111
rect 569408 445800 569460 445806
rect 569408 445742 569460 445748
rect 569408 431588 569460 431594
rect 569408 431530 569460 431536
rect 569420 431497 569448 431530
rect 569406 431488 569462 431497
rect 569406 431423 569462 431432
rect 569316 365696 569368 365702
rect 569316 365638 569368 365644
rect 569314 321872 569370 321881
rect 569314 321807 569370 321816
rect 569328 321638 569356 321807
rect 569316 321632 569368 321638
rect 569316 321574 569368 321580
rect 569314 266520 569370 266529
rect 569314 266455 569370 266464
rect 569328 266422 569356 266455
rect 569316 266416 569368 266422
rect 569316 266358 569368 266364
rect 569314 258632 569370 258641
rect 569314 258567 569370 258576
rect 569328 258534 569356 258567
rect 569316 258528 569368 258534
rect 569316 258470 569368 258476
rect 569590 242856 569646 242865
rect 569590 242791 569646 242800
rect 569314 235104 569370 235113
rect 569314 235039 569370 235048
rect 569328 71194 569356 235039
rect 569406 219872 569462 219881
rect 569406 219807 569462 219816
rect 569420 219774 569448 219807
rect 569408 219768 569460 219774
rect 569408 219710 569460 219716
rect 569406 204096 569462 204105
rect 569406 204031 569462 204040
rect 569316 71188 569368 71194
rect 569316 71130 569368 71136
rect 569314 71088 569370 71097
rect 569314 71023 569370 71032
rect 569328 68406 569356 71023
rect 569420 69018 569448 204031
rect 569498 149152 569554 149161
rect 569498 149087 569554 149096
rect 569408 69012 569460 69018
rect 569408 68954 569460 68960
rect 569316 68400 569368 68406
rect 569316 68342 569368 68348
rect 569512 64190 569540 149087
rect 569604 69290 569632 242791
rect 569972 126857 570000 683130
rect 570064 158137 570092 700266
rect 570236 566500 570288 566506
rect 570236 566442 570288 566448
rect 570142 540560 570198 540569
rect 570142 540495 570198 540504
rect 570050 158128 570106 158137
rect 570050 158063 570106 158072
rect 570050 133920 570106 133929
rect 570050 133855 570106 133864
rect 569958 126848 570014 126857
rect 569958 126783 570014 126792
rect 569682 117872 569738 117881
rect 569682 117807 569738 117816
rect 569592 69284 569644 69290
rect 569592 69226 569644 69232
rect 569696 68882 569724 117807
rect 569958 87408 570014 87417
rect 569958 87343 570014 87352
rect 569776 80096 569828 80102
rect 569776 80038 569828 80044
rect 569684 68876 569736 68882
rect 569684 68818 569736 68824
rect 569500 64184 569552 64190
rect 569500 64126 569552 64132
rect 569788 3670 569816 80038
rect 569868 71188 569920 71194
rect 569868 71130 569920 71136
rect 569880 67046 569908 71130
rect 569972 68814 570000 87343
rect 569960 68808 570012 68814
rect 569960 68750 570012 68756
rect 570064 68542 570092 133855
rect 570052 68536 570104 68542
rect 570052 68478 570104 68484
rect 570156 68134 570184 540495
rect 570248 165209 570276 566442
rect 570340 517177 570368 700538
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 576216 683188 576268 683194
rect 576216 683130 576268 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 573364 670744 573416 670750
rect 573364 670686 573416 670692
rect 570420 632120 570472 632126
rect 570420 632062 570472 632068
rect 570326 517168 570382 517177
rect 570326 517103 570382 517112
rect 570326 462496 570382 462505
rect 570326 462431 570382 462440
rect 570234 165200 570290 165209
rect 570234 165135 570290 165144
rect 570234 95024 570290 95033
rect 570234 94959 570290 94968
rect 570248 68610 570276 94959
rect 570340 70038 570368 462431
rect 570432 423337 570460 632062
rect 571248 567316 571300 567322
rect 571248 567258 571300 567264
rect 570604 567248 570656 567254
rect 570604 567190 570656 567196
rect 570616 458182 570644 567190
rect 571260 564398 571288 567258
rect 571248 564392 571300 564398
rect 571248 564334 571300 564340
rect 571338 556064 571394 556073
rect 571338 555999 571394 556008
rect 571352 554810 571380 555999
rect 571340 554804 571392 554810
rect 571340 554746 571392 554752
rect 571706 532672 571762 532681
rect 571706 532607 571762 532616
rect 571430 485888 571486 485897
rect 571430 485823 571486 485832
rect 571338 478000 571394 478009
rect 571338 477935 571394 477944
rect 571352 477698 571380 477935
rect 571340 477692 571392 477698
rect 571340 477634 571392 477640
rect 570604 458176 570656 458182
rect 570604 458118 570656 458124
rect 570418 423328 570474 423337
rect 570418 423263 570474 423272
rect 570418 407552 570474 407561
rect 570418 407487 570474 407496
rect 570328 70032 570380 70038
rect 570328 69974 570380 69980
rect 570432 68950 570460 407487
rect 570510 399936 570566 399945
rect 570510 399871 570566 399880
rect 570524 69970 570552 399871
rect 571338 306096 571394 306105
rect 571338 306031 571394 306040
rect 571352 305658 571380 306031
rect 571340 305652 571392 305658
rect 571340 305594 571392 305600
rect 570602 274816 570658 274825
rect 570602 274751 570658 274760
rect 570616 70106 570644 274751
rect 570694 212256 570750 212265
rect 570694 212191 570750 212200
rect 570604 70100 570656 70106
rect 570604 70042 570656 70048
rect 570512 69964 570564 69970
rect 570512 69906 570564 69912
rect 570420 68944 570472 68950
rect 570420 68886 570472 68892
rect 570236 68604 570288 68610
rect 570236 68546 570288 68552
rect 570708 68202 570736 212191
rect 570878 196480 570934 196489
rect 570878 196415 570934 196424
rect 570788 140820 570840 140826
rect 570788 140762 570840 140768
rect 570696 68196 570748 68202
rect 570696 68138 570748 68144
rect 570144 68128 570196 68134
rect 570144 68070 570196 68076
rect 569868 67040 569920 67046
rect 569868 66982 569920 66988
rect 569776 3664 569828 3670
rect 569776 3606 569828 3612
rect 570800 3534 570828 140762
rect 570892 66910 570920 196415
rect 570970 188864 571026 188873
rect 570970 188799 571026 188808
rect 570984 69902 571012 188799
rect 571338 79248 571394 79257
rect 571338 79183 571394 79192
rect 570972 69896 571024 69902
rect 570972 69838 571024 69844
rect 571352 69698 571380 79183
rect 571340 69692 571392 69698
rect 571340 69634 571392 69640
rect 571444 69630 571472 485823
rect 571522 470112 571578 470121
rect 571522 470047 571578 470056
rect 571536 80102 571564 470047
rect 571614 415440 571670 415449
rect 571614 415375 571670 415384
rect 571524 80096 571576 80102
rect 571524 80038 571576 80044
rect 571432 69624 571484 69630
rect 571432 69566 571484 69572
rect 570880 66904 570932 66910
rect 570880 66846 570932 66852
rect 571628 65890 571656 415375
rect 571720 390590 571748 532607
rect 571982 524784 572038 524793
rect 571982 524719 572038 524728
rect 571996 511970 572024 524719
rect 571984 511964 572036 511970
rect 571984 511906 572036 511912
rect 572442 509280 572498 509289
rect 572442 509215 572498 509224
rect 571708 390584 571760 390590
rect 571708 390526 571760 390532
rect 571798 384160 571854 384169
rect 571798 384095 571854 384104
rect 571706 141808 571762 141817
rect 571706 141743 571762 141752
rect 571720 132494 571748 141743
rect 571812 140826 571840 384095
rect 572076 345024 572128 345030
rect 572074 344992 572076 345001
rect 572128 344992 572130 345001
rect 572074 344927 572130 344936
rect 571890 298208 571946 298217
rect 571890 298143 571946 298152
rect 571800 140820 571852 140826
rect 571800 140762 571852 140768
rect 571720 132466 571840 132494
rect 571812 68270 571840 132466
rect 571904 69222 571932 298143
rect 571982 282704 572038 282713
rect 571982 282639 572038 282648
rect 571996 69834 572024 282639
rect 572074 251424 572130 251433
rect 572074 251359 572130 251368
rect 571984 69828 572036 69834
rect 571984 69770 572036 69776
rect 572088 69766 572116 251359
rect 572166 227760 572222 227769
rect 572166 227695 572222 227704
rect 572076 69760 572128 69766
rect 572076 69702 572128 69708
rect 571892 69216 571944 69222
rect 571892 69158 571944 69164
rect 572180 68338 572208 227695
rect 572258 110528 572314 110537
rect 572258 110463 572314 110472
rect 572272 69426 572300 110463
rect 572350 102912 572406 102921
rect 572350 102847 572406 102856
rect 572260 69420 572312 69426
rect 572260 69362 572312 69368
rect 572168 68332 572220 68338
rect 572168 68274 572220 68280
rect 571800 68264 571852 68270
rect 571800 68206 571852 68212
rect 572364 67182 572392 102847
rect 572456 68678 572484 509215
rect 572626 454608 572682 454617
rect 572682 454566 572760 454594
rect 572626 454543 572682 454552
rect 572534 392048 572590 392057
rect 572534 391983 572590 391992
rect 572548 68746 572576 391983
rect 572628 329588 572680 329594
rect 572628 329530 572680 329536
rect 572640 329497 572668 329530
rect 572626 329488 572682 329497
rect 572626 329423 572682 329432
rect 572536 68740 572588 68746
rect 572536 68682 572588 68688
rect 572444 68672 572496 68678
rect 572444 68614 572496 68620
rect 572352 67176 572404 67182
rect 572352 67118 572404 67124
rect 571616 65884 571668 65890
rect 571616 65826 571668 65832
rect 572732 62830 572760 454566
rect 572810 360768 572866 360777
rect 572810 360703 572866 360712
rect 572720 62824 572772 62830
rect 572720 62766 572772 62772
rect 572824 6186 572852 360703
rect 572902 352880 572958 352889
rect 572902 352815 572958 352824
rect 572916 6322 572944 352815
rect 572996 305652 573048 305658
rect 572996 305594 573048 305600
rect 572904 6316 572956 6322
rect 572904 6258 572956 6264
rect 572812 6180 572864 6186
rect 572812 6122 572864 6128
rect 573008 4894 573036 305594
rect 573376 66706 573404 670686
rect 574744 576904 574796 576910
rect 574744 576846 574796 576852
rect 573456 568268 573508 568274
rect 573456 568210 573508 568216
rect 573364 66700 573416 66706
rect 573364 66642 573416 66648
rect 573468 60722 573496 568210
rect 573548 567928 573600 567934
rect 573548 567870 573600 567876
rect 573560 126954 573588 567870
rect 573732 554804 573784 554810
rect 573732 554746 573784 554752
rect 573640 477692 573692 477698
rect 573640 477634 573692 477640
rect 573652 139398 573680 477634
rect 573744 405686 573772 554746
rect 573732 405680 573784 405686
rect 573732 405622 573784 405628
rect 573640 139392 573692 139398
rect 573640 139334 573692 139340
rect 573548 126948 573600 126954
rect 573548 126890 573600 126896
rect 574756 66094 574784 576846
rect 574928 567656 574980 567662
rect 574928 567598 574980 567604
rect 574836 567520 574888 567526
rect 574836 567462 574888 567468
rect 574848 167006 574876 567462
rect 574940 245614 574968 567598
rect 576124 567452 576176 567458
rect 576124 567394 576176 567400
rect 575020 418192 575072 418198
rect 575020 418134 575072 418140
rect 575032 345030 575060 418134
rect 575020 345024 575072 345030
rect 575020 344966 575072 344972
rect 575020 258120 575072 258126
rect 575020 258062 575072 258068
rect 574928 245608 574980 245614
rect 574928 245550 574980 245556
rect 574928 218068 574980 218074
rect 574928 218010 574980 218016
rect 574836 167000 574888 167006
rect 574836 166942 574888 166948
rect 574940 67250 574968 218010
rect 574928 67244 574980 67250
rect 574928 67186 574980 67192
rect 575032 66230 575060 258062
rect 576136 100706 576164 567394
rect 576228 329594 576256 683130
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 576308 568132 576360 568138
rect 576308 568074 576360 568080
rect 576216 329588 576268 329594
rect 576216 329530 576268 329536
rect 576320 299470 576348 568074
rect 580264 568064 580316 568070
rect 580264 568006 580316 568012
rect 577504 567996 577556 568002
rect 577504 567938 577556 567944
rect 576308 299464 576360 299470
rect 576308 299406 576360 299412
rect 577516 179382 577544 567938
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580276 524521 580304 568006
rect 580356 567792 580408 567798
rect 580356 567734 580408 567740
rect 580262 524512 580318 524521
rect 580262 524447 580318 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580262 471472 580318 471481
rect 580262 471407 580318 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 579988 365696 580040 365702
rect 579988 365638 580040 365644
rect 580000 365129 580028 365638
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579632 258126 579660 258839
rect 579620 258120 579672 258126
rect 579620 258062 579672 258068
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 577504 179376 577556 179382
rect 577504 179318 577556 179324
rect 579896 179376 579948 179382
rect 579896 179318 579948 179324
rect 579908 179217 579936 179318
rect 579894 179208 579950 179217
rect 579894 179143 579950 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 576124 100700 576176 100706
rect 576124 100642 576176 100648
rect 579712 100700 579764 100706
rect 579712 100642 579764 100648
rect 579724 99521 579752 100642
rect 579710 99512 579766 99521
rect 579710 99447 579766 99456
rect 580276 69494 580304 471407
rect 580368 351937 580396 567734
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580354 312080 580410 312089
rect 580354 312015 580410 312024
rect 580264 69488 580316 69494
rect 580264 69430 580316 69436
rect 580264 66972 580316 66978
rect 580264 66914 580316 66920
rect 575020 66224 575072 66230
rect 575020 66166 575072 66172
rect 574744 66088 574796 66094
rect 574744 66030 574796 66036
rect 573456 60716 573508 60722
rect 573456 60658 573508 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 580276 6633 580304 66914
rect 580368 66842 580396 312015
rect 580446 205728 580502 205737
rect 580446 205663 580502 205672
rect 580356 66836 580408 66842
rect 580356 66778 580408 66784
rect 580460 66774 580488 205663
rect 580538 86184 580594 86193
rect 580538 86119 580594 86128
rect 580552 69562 580580 86119
rect 580540 69556 580592 69562
rect 580540 69498 580592 69504
rect 580448 66768 580500 66774
rect 580448 66710 580500 66716
rect 580356 55888 580408 55894
rect 580356 55830 580408 55836
rect 580368 46345 580396 55830
rect 580354 46336 580410 46345
rect 580354 46271 580410 46280
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 572996 4888 573048 4894
rect 572996 4830 573048 4836
rect 570788 3528 570840 3534
rect 570788 3470 570840 3476
rect 569224 3460 569276 3466
rect 569224 3402 569276 3408
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 671200 2834 671256
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3514 619112 3570 619168
rect 2778 579964 2834 580000
rect 2778 579944 2780 579964
rect 2780 579944 2832 579964
rect 2832 579944 2834 579964
rect 3514 566888 3570 566944
rect 3514 527856 3570 527912
rect 3422 514800 3478 514856
rect 2778 475632 2834 475688
rect 3422 462576 3478 462632
rect 2778 423564 2834 423600
rect 2778 423544 2780 423564
rect 2780 423544 2832 423564
rect 2832 423544 2834 423564
rect 3330 410488 3386 410544
rect 3330 358400 3386 358456
rect 3238 214920 3294 214976
rect 2778 149776 2834 149832
rect 3330 97552 3386 97608
rect 3606 371320 3662 371376
rect 3514 319232 3570 319288
rect 3514 306176 3570 306232
rect 3790 267144 3846 267200
rect 3698 162832 3754 162888
rect 3606 110608 3662 110664
rect 4066 254088 4122 254144
rect 3974 201864 4030 201920
rect 3882 71576 3938 71632
rect 3054 58520 3110 58576
rect 3698 32408 3754 32464
rect 3422 19352 3478 19408
rect 67638 560360 67694 560416
rect 68742 552472 68798 552528
rect 67546 544856 67602 544912
rect 67454 529080 67510 529136
rect 67362 521192 67418 521248
rect 67270 505688 67326 505744
rect 67178 435240 67234 435296
rect 67086 419736 67142 419792
rect 66994 224168 67050 224224
rect 66902 185272 66958 185328
rect 67638 536968 67694 537024
rect 68742 513576 68798 513632
rect 68650 497800 68706 497856
rect 68374 482296 68430 482352
rect 68282 474408 68338 474464
rect 67914 427352 67970 427408
rect 67638 411848 67694 411904
rect 68006 403960 68062 404016
rect 67638 396344 67694 396400
rect 67638 372680 67694 372736
rect 67638 365064 67694 365120
rect 67822 357176 67878 357232
rect 67638 349288 67694 349344
rect 67638 325896 67694 325952
rect 67822 302504 67878 302560
rect 67822 286728 67878 286784
rect 68190 278840 68246 278896
rect 67638 271224 67694 271280
rect 68282 263336 68338 263392
rect 68190 255448 68246 255504
rect 67638 239944 67694 240000
rect 67638 232056 67694 232112
rect 67638 208664 67694 208720
rect 67730 200776 67786 200832
rect 67638 177384 67694 177440
rect 67638 161608 67694 161664
rect 67638 138216 67694 138272
rect 67638 130328 67694 130384
rect 67638 99048 67694 99104
rect 67638 91432 67694 91488
rect 68098 192888 68154 192944
rect 68006 153992 68062 154048
rect 67914 146104 67970 146160
rect 67822 114824 67878 114880
rect 68098 122712 68154 122768
rect 68558 466520 68614 466576
rect 68466 443128 68522 443184
rect 68374 247560 68430 247616
rect 68374 83544 68430 83600
rect 68650 451016 68706 451072
rect 69018 388456 69074 388512
rect 69202 318008 69258 318064
rect 69110 310120 69166 310176
rect 69294 294616 69350 294672
rect 105450 699760 105506 699816
rect 235170 699760 235226 699816
rect 249982 571240 250038 571296
rect 176014 570968 176070 571024
rect 178130 568520 178186 568576
rect 302790 571104 302846 571160
rect 292302 570832 292358 570888
rect 286966 570696 287022 570752
rect 297454 570560 297510 570616
rect 392766 570968 392822 571024
rect 349986 570832 350042 570888
rect 376942 570696 376998 570752
rect 349986 570560 350042 570616
rect 382094 570424 382150 570480
rect 413926 570288 413982 570344
rect 403254 570152 403310 570208
rect 429842 699760 429898 699816
rect 519542 570560 519598 570616
rect 524878 570016 524934 570072
rect 546038 570152 546094 570208
rect 86406 567296 86462 567352
rect 102046 567296 102102 567352
rect 128634 567296 128690 567352
rect 133510 567296 133566 567352
rect 144550 567296 144606 567352
rect 155222 567296 155278 567352
rect 170954 567296 171010 567352
rect 212722 567296 212778 567352
rect 228546 567296 228602 567352
rect 244370 567296 244426 567352
rect 270866 567296 270922 567352
rect 281446 567296 281502 567352
rect 329010 567296 329066 567352
rect 339590 567296 339646 567352
rect 345294 567296 345350 567352
rect 387154 567296 387210 567352
rect 440054 567296 440110 567352
rect 461122 567296 461178 567352
rect 482282 567296 482338 567352
rect 540426 567296 540482 567352
rect 551098 567296 551154 567352
rect 92754 3440 92810 3496
rect 97446 3440 97502 3496
rect 109314 5208 109370 5264
rect 108118 4936 108174 4992
rect 106922 3576 106978 3632
rect 105726 3304 105782 3360
rect 110510 3440 110566 3496
rect 118790 4800 118846 4856
rect 117594 3576 117650 3632
rect 130566 3712 130622 3768
rect 135258 5072 135314 5128
rect 140042 3712 140098 3768
rect 145930 3712 145986 3768
rect 150622 6704 150678 6760
rect 153014 3712 153070 3768
rect 156602 3712 156658 3768
rect 161294 5888 161350 5944
rect 160098 3712 160154 3768
rect 166078 5480 166134 5536
rect 164882 3712 164938 3768
rect 180982 67224 181038 67280
rect 168378 5072 168434 5128
rect 170770 4936 170826 4992
rect 180246 6160 180302 6216
rect 183742 6024 183798 6080
rect 195610 6296 195666 6352
rect 200302 6568 200358 6624
rect 201498 5344 201554 5400
rect 203890 5208 203946 5264
rect 205086 3576 205142 3632
rect 210974 3576 211030 3632
rect 223302 67496 223358 67552
rect 220450 3576 220506 3632
rect 226338 6840 226394 6896
rect 227534 3576 227590 3632
rect 233422 6432 233478 6488
rect 237010 6432 237066 6488
rect 238114 5072 238170 5128
rect 307942 67360 307998 67416
rect 569406 564304 569462 564360
rect 569406 548140 569462 548176
rect 569406 548120 569408 548140
rect 569408 548120 569460 548140
rect 569460 548120 569462 548140
rect 569406 500792 569462 500848
rect 569406 493992 569462 494048
rect 569406 446120 569462 446176
rect 569406 431432 569462 431488
rect 569314 321816 569370 321872
rect 569314 266464 569370 266520
rect 569314 258576 569370 258632
rect 569590 242800 569646 242856
rect 569314 235048 569370 235104
rect 569406 219816 569462 219872
rect 569406 204040 569462 204096
rect 569314 71032 569370 71088
rect 569498 149096 569554 149152
rect 570142 540504 570198 540560
rect 570050 158072 570106 158128
rect 570050 133864 570106 133920
rect 569958 126792 570014 126848
rect 569682 117816 569738 117872
rect 569958 87352 570014 87408
rect 580170 683848 580226 683904
rect 570326 517112 570382 517168
rect 570326 462440 570382 462496
rect 570234 165144 570290 165200
rect 570234 94968 570290 95024
rect 571338 556008 571394 556064
rect 571706 532616 571762 532672
rect 571430 485832 571486 485888
rect 571338 477944 571394 478000
rect 570418 423272 570474 423328
rect 570418 407496 570474 407552
rect 570510 399880 570566 399936
rect 571338 306040 571394 306096
rect 570602 274760 570658 274816
rect 570694 212200 570750 212256
rect 570878 196424 570934 196480
rect 570970 188808 571026 188864
rect 571338 79192 571394 79248
rect 571522 470056 571578 470112
rect 571614 415384 571670 415440
rect 571982 524728 572038 524784
rect 572442 509224 572498 509280
rect 571798 384104 571854 384160
rect 571706 141752 571762 141808
rect 572074 344972 572076 344992
rect 572076 344972 572128 344992
rect 572128 344972 572130 344992
rect 572074 344936 572130 344972
rect 571890 298152 571946 298208
rect 571982 282648 572038 282704
rect 572074 251368 572130 251424
rect 572166 227704 572222 227760
rect 572258 110472 572314 110528
rect 572350 102856 572406 102912
rect 572626 454552 572682 454608
rect 572534 391992 572590 392048
rect 572626 329432 572682 329488
rect 572810 360712 572866 360768
rect 572902 352824 572958 352880
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580170 577632 580226 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580262 524456 580318 524512
rect 580170 511264 580226 511320
rect 580262 471416 580318 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 579986 365064 580042 365120
rect 580170 298696 580226 298752
rect 579618 258848 579674 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 219000 580226 219056
rect 579894 179152 579950 179208
rect 580170 165824 580226 165880
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579618 125976 579674 126032
rect 579710 99456 579766 99512
rect 580354 351872 580410 351928
rect 580354 312024 580410 312080
rect 580170 59608 580226 59664
rect 580170 19760 580226 19816
rect 580446 205672 580502 205728
rect 580538 86128 580594 86184
rect 580354 46280 580410 46336
rect 580262 6568 580318 6624
<< metal3 >>
rect 105445 699818 105511 699821
rect 106774 699818 106780 699820
rect 105445 699816 106780 699818
rect 105445 699760 105450 699816
rect 105506 699760 106780 699816
rect 105445 699758 106780 699760
rect 105445 699755 105511 699758
rect 106774 699756 106780 699758
rect 106844 699756 106850 699820
rect 234654 699756 234660 699820
rect 234724 699818 234730 699820
rect 235165 699818 235231 699821
rect 234724 699816 235231 699818
rect 234724 699760 235170 699816
rect 235226 699760 235231 699816
rect 234724 699758 235231 699760
rect 234724 699756 234730 699758
rect 235165 699755 235231 699758
rect 429142 699756 429148 699820
rect 429212 699818 429218 699820
rect 429837 699818 429903 699821
rect 429212 699816 429903 699818
rect 429212 699760 429842 699816
rect 429898 699760 429903 699816
rect 429212 699758 429903 699760
rect 429212 699756 429218 699758
rect 429837 699755 429903 699758
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 152958 571236 152964 571300
rect 153028 571298 153034 571300
rect 249977 571298 250043 571301
rect 153028 571296 250043 571298
rect 153028 571240 249982 571296
rect 250038 571240 250043 571296
rect 153028 571238 250043 571240
rect 153028 571236 153034 571238
rect 249977 571235 250043 571238
rect 175774 571100 175780 571164
rect 175844 571162 175850 571164
rect 302785 571162 302851 571165
rect 175844 571160 302851 571162
rect 175844 571104 302790 571160
rect 302846 571104 302851 571160
rect 175844 571102 302851 571104
rect 175844 571100 175850 571102
rect 302785 571099 302851 571102
rect 156638 570964 156644 571028
rect 156708 571026 156714 571028
rect 176009 571026 176075 571029
rect 156708 571024 176075 571026
rect 156708 570968 176014 571024
rect 176070 570968 176075 571024
rect 156708 570966 176075 570968
rect 156708 570964 156714 570966
rect 176009 570963 176075 570966
rect 227478 570964 227484 571028
rect 227548 571026 227554 571028
rect 392761 571026 392827 571029
rect 227548 571024 392827 571026
rect 227548 570968 392766 571024
rect 392822 570968 392827 571024
rect 227548 570966 392827 570968
rect 227548 570964 227554 570966
rect 392761 570963 392827 570966
rect 111558 570828 111564 570892
rect 111628 570890 111634 570892
rect 292297 570890 292363 570893
rect 111628 570888 292363 570890
rect 111628 570832 292302 570888
rect 292358 570832 292363 570888
rect 111628 570830 292363 570832
rect 111628 570828 111634 570830
rect 292297 570827 292363 570830
rect 346894 570828 346900 570892
rect 346964 570890 346970 570892
rect 349981 570890 350047 570893
rect 346964 570888 350047 570890
rect 346964 570832 349986 570888
rect 350042 570832 350047 570888
rect 346964 570830 350047 570832
rect 346964 570828 346970 570830
rect 349981 570827 350047 570830
rect 93710 570692 93716 570756
rect 93780 570754 93786 570756
rect 286961 570754 287027 570757
rect 93780 570752 287027 570754
rect 93780 570696 286966 570752
rect 287022 570696 287027 570752
rect 93780 570694 287027 570696
rect 93780 570692 93786 570694
rect 286961 570691 287027 570694
rect 348366 570692 348372 570756
rect 348436 570754 348442 570756
rect 376937 570754 377003 570757
rect 348436 570752 377003 570754
rect 348436 570696 376942 570752
rect 376998 570696 377003 570752
rect 348436 570694 377003 570696
rect 348436 570692 348442 570694
rect 376937 570691 377003 570694
rect 97758 570556 97764 570620
rect 97828 570618 97834 570620
rect 297449 570618 297515 570621
rect 349981 570618 350047 570621
rect 519537 570618 519603 570621
rect 97828 570616 297515 570618
rect 97828 570560 297454 570616
rect 297510 570560 297515 570616
rect 97828 570558 297515 570560
rect 97828 570556 97834 570558
rect 297449 570555 297515 570558
rect 315990 570558 349906 570618
rect 168966 570420 168972 570484
rect 169036 570482 169042 570484
rect 315990 570482 316050 570558
rect 349846 570482 349906 570558
rect 349981 570616 519603 570618
rect 349981 570560 349986 570616
rect 350042 570560 519542 570616
rect 519598 570560 519603 570616
rect 349981 570558 519603 570560
rect 349981 570555 350047 570558
rect 519537 570555 519603 570558
rect 382089 570482 382155 570485
rect 169036 570422 316050 570482
rect 335310 570422 349722 570482
rect 349846 570480 382155 570482
rect 349846 570424 382094 570480
rect 382150 570424 382155 570480
rect 349846 570422 382155 570424
rect 169036 570420 169042 570422
rect 161238 570284 161244 570348
rect 161308 570346 161314 570348
rect 335310 570346 335370 570422
rect 349662 570346 349722 570422
rect 382089 570419 382155 570422
rect 413921 570346 413987 570349
rect 161308 570286 335370 570346
rect 344970 570286 349538 570346
rect 349662 570344 413987 570346
rect 349662 570288 413926 570344
rect 413982 570288 413987 570344
rect 349662 570286 413987 570288
rect 161308 570284 161314 570286
rect 145598 570148 145604 570212
rect 145668 570210 145674 570212
rect 344970 570210 345030 570286
rect 145668 570150 345030 570210
rect 349478 570210 349538 570286
rect 413921 570283 413987 570286
rect 403249 570210 403315 570213
rect 349478 570208 403315 570210
rect 349478 570152 403254 570208
rect 403310 570152 403315 570208
rect 349478 570150 403315 570152
rect 145668 570148 145674 570150
rect 403249 570147 403315 570150
rect 403566 570148 403572 570212
rect 403636 570210 403642 570212
rect 546033 570210 546099 570213
rect 403636 570208 546099 570210
rect 403636 570152 546038 570208
rect 546094 570152 546099 570208
rect 403636 570150 546099 570152
rect 403636 570148 403642 570150
rect 546033 570147 546099 570150
rect 220670 570012 220676 570076
rect 220740 570074 220746 570076
rect 524873 570074 524939 570077
rect 220740 570072 524939 570074
rect 220740 570016 524878 570072
rect 524934 570016 524939 570072
rect 220740 570014 524939 570016
rect 220740 570012 220746 570014
rect 524873 570011 524939 570014
rect 177982 568516 177988 568580
rect 178052 568578 178058 568580
rect 178125 568578 178191 568581
rect 178052 568576 178191 568578
rect 178052 568520 178130 568576
rect 178186 568520 178191 568576
rect 178052 568518 178191 568520
rect 178052 568516 178058 568518
rect 178125 568515 178191 568518
rect 86401 567354 86467 567357
rect 102041 567356 102107 567357
rect 86718 567354 86724 567356
rect 86401 567352 86724 567354
rect 86401 567296 86406 567352
rect 86462 567296 86724 567352
rect 86401 567294 86724 567296
rect 86401 567291 86467 567294
rect 86718 567292 86724 567294
rect 86788 567292 86794 567356
rect 101990 567354 101996 567356
rect 101950 567294 101996 567354
rect 102060 567352 102107 567356
rect 102102 567296 102107 567352
rect 101990 567292 101996 567294
rect 102060 567292 102107 567296
rect 102041 567291 102107 567292
rect 128629 567354 128695 567357
rect 133505 567354 133571 567357
rect 133638 567354 133644 567356
rect 128629 567352 128738 567354
rect 128629 567296 128634 567352
rect 128690 567296 128738 567352
rect 128629 567291 128738 567296
rect 133505 567352 133644 567354
rect 133505 567296 133510 567352
rect 133566 567296 133644 567352
rect 133505 567294 133644 567296
rect 133505 567291 133571 567294
rect 133638 567292 133644 567294
rect 133708 567292 133714 567356
rect 144545 567354 144611 567357
rect 144678 567354 144684 567356
rect 144545 567352 144684 567354
rect 144545 567296 144550 567352
rect 144606 567296 144684 567352
rect 144545 567294 144684 567296
rect 144545 567291 144611 567294
rect 144678 567292 144684 567294
rect 144748 567292 144754 567356
rect 155217 567354 155283 567357
rect 170949 567356 171015 567357
rect 155718 567354 155724 567356
rect 155217 567352 155724 567354
rect 155217 567296 155222 567352
rect 155278 567296 155724 567352
rect 155217 567294 155724 567296
rect 155217 567291 155283 567294
rect 155718 567292 155724 567294
rect 155788 567292 155794 567356
rect 170949 567352 170996 567356
rect 171060 567354 171066 567356
rect 170949 567296 170954 567352
rect 170949 567292 170996 567296
rect 171060 567294 171106 567354
rect 171060 567292 171066 567294
rect 210366 567292 210372 567356
rect 210436 567354 210442 567356
rect 212717 567354 212783 567357
rect 228541 567354 228607 567357
rect 210436 567352 212783 567354
rect 210436 567296 212722 567352
rect 212778 567296 212783 567352
rect 210436 567294 212783 567296
rect 210436 567292 210442 567294
rect 170949 567291 171015 567292
rect 212717 567291 212783 567294
rect 219390 567352 228607 567354
rect 219390 567296 228546 567352
rect 228602 567296 228607 567352
rect 219390 567294 228607 567296
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 128678 566674 128738 567291
rect 214414 567156 214420 567220
rect 214484 567218 214490 567220
rect 219390 567218 219450 567294
rect 228541 567291 228607 567294
rect 244222 567292 244228 567356
rect 244292 567354 244298 567356
rect 244365 567354 244431 567357
rect 244292 567352 244431 567354
rect 244292 567296 244370 567352
rect 244426 567296 244431 567352
rect 244292 567294 244431 567296
rect 244292 567292 244298 567294
rect 244365 567291 244431 567294
rect 270534 567292 270540 567356
rect 270604 567354 270610 567356
rect 270861 567354 270927 567357
rect 270604 567352 270927 567354
rect 270604 567296 270866 567352
rect 270922 567296 270927 567352
rect 270604 567294 270927 567296
rect 270604 567292 270610 567294
rect 270861 567291 270927 567294
rect 281441 567354 281507 567357
rect 281574 567354 281580 567356
rect 281441 567352 281580 567354
rect 281441 567296 281446 567352
rect 281502 567296 281580 567352
rect 281441 567294 281580 567296
rect 281441 567291 281507 567294
rect 281574 567292 281580 567294
rect 281644 567292 281650 567356
rect 328494 567292 328500 567356
rect 328564 567354 328570 567356
rect 329005 567354 329071 567357
rect 339585 567354 339651 567357
rect 328564 567352 329071 567354
rect 328564 567296 329010 567352
rect 329066 567296 329071 567352
rect 328564 567294 329071 567296
rect 328564 567292 328570 567294
rect 329005 567291 329071 567294
rect 339542 567352 339651 567354
rect 339542 567296 339590 567352
rect 339646 567296 339651 567352
rect 339542 567291 339651 567296
rect 345054 567292 345060 567356
rect 345124 567354 345130 567356
rect 345289 567354 345355 567357
rect 345124 567352 345355 567354
rect 345124 567296 345294 567352
rect 345350 567296 345355 567352
rect 345124 567294 345355 567296
rect 345124 567292 345130 567294
rect 345289 567291 345355 567294
rect 386454 567292 386460 567356
rect 386524 567354 386530 567356
rect 387149 567354 387215 567357
rect 386524 567352 387215 567354
rect 386524 567296 387154 567352
rect 387210 567296 387215 567352
rect 386524 567294 387215 567296
rect 386524 567292 386530 567294
rect 387149 567291 387215 567294
rect 440049 567354 440115 567357
rect 440182 567354 440188 567356
rect 440049 567352 440188 567354
rect 440049 567296 440054 567352
rect 440110 567296 440188 567352
rect 440049 567294 440188 567296
rect 440049 567291 440115 567294
rect 440182 567292 440188 567294
rect 440252 567292 440258 567356
rect 460974 567292 460980 567356
rect 461044 567354 461050 567356
rect 461117 567354 461183 567357
rect 461044 567352 461183 567354
rect 461044 567296 461122 567352
rect 461178 567296 461183 567352
rect 461044 567294 461183 567296
rect 461044 567292 461050 567294
rect 461117 567291 461183 567294
rect 481766 567292 481772 567356
rect 481836 567354 481842 567356
rect 482277 567354 482343 567357
rect 481836 567352 482343 567354
rect 481836 567296 482282 567352
rect 482338 567296 482343 567352
rect 481836 567294 482343 567296
rect 481836 567292 481842 567294
rect 482277 567291 482343 567294
rect 539542 567292 539548 567356
rect 539612 567354 539618 567356
rect 540421 567354 540487 567357
rect 539612 567352 540487 567354
rect 539612 567296 540426 567352
rect 540482 567296 540487 567352
rect 539612 567294 540487 567296
rect 539612 567292 539618 567294
rect 540421 567291 540487 567294
rect 550766 567292 550772 567356
rect 550836 567354 550842 567356
rect 551093 567354 551159 567357
rect 550836 567352 551159 567354
rect 550836 567296 551098 567352
rect 551154 567296 551159 567352
rect 550836 567294 551159 567296
rect 550836 567292 550842 567294
rect 551093 567291 551159 567294
rect 214484 567158 219450 567218
rect 214484 567156 214490 567158
rect 164550 566674 164556 566676
rect 128678 566614 164556 566674
rect 164550 566612 164556 566614
rect 164620 566612 164626 566676
rect 130878 566476 130884 566540
rect 130948 566538 130954 566540
rect 328494 566538 328500 566540
rect 130948 566478 328500 566538
rect 130948 566476 130954 566478
rect 328494 566476 328500 566478
rect 328564 566476 328570 566540
rect 140630 566340 140636 566404
rect 140700 566402 140706 566404
rect 339542 566402 339602 567291
rect 140700 566342 339602 566402
rect 140700 566340 140706 566342
rect 205398 565932 205404 565996
rect 205468 565994 205474 565996
rect 210366 565994 210372 565996
rect 205468 565934 210372 565994
rect 205468 565932 205474 565934
rect 210366 565932 210372 565934
rect 210436 565932 210442 565996
rect 569401 564362 569467 564365
rect 569358 564360 569467 564362
rect 569358 564304 569406 564360
rect 569462 564304 569467 564360
rect 569358 564299 569467 564304
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 569358 563924 569418 564299
rect 583520 564212 584960 564302
rect 67633 560418 67699 560421
rect 67633 560416 70012 560418
rect 67633 560360 67638 560416
rect 67694 560360 70012 560416
rect 67633 560358 70012 560360
rect 67633 560355 67699 560358
rect 571333 556066 571399 556069
rect 569940 556064 571399 556066
rect 569940 556008 571338 556064
rect 571394 556008 571399 556064
rect 569940 556006 571399 556008
rect 571333 556003 571399 556006
rect -960 553740 480 553980
rect 68737 552530 68803 552533
rect 68737 552528 70012 552530
rect 68737 552472 68742 552528
rect 68798 552472 70012 552528
rect 68737 552470 70012 552472
rect 68737 552467 68803 552470
rect 583520 551020 584960 551260
rect 569358 548181 569418 548420
rect 569358 548176 569467 548181
rect 569358 548120 569406 548176
rect 569462 548120 569467 548176
rect 569358 548118 569467 548120
rect 569401 548115 569467 548118
rect 67541 544914 67607 544917
rect 67541 544912 70012 544914
rect 67541 544856 67546 544912
rect 67602 544856 70012 544912
rect 67541 544854 70012 544856
rect 67541 544851 67607 544854
rect -960 540684 480 540924
rect 570137 540562 570203 540565
rect 569940 540560 570203 540562
rect 569940 540504 570142 540560
rect 570198 540504 570203 540560
rect 569940 540502 570203 540504
rect 570137 540499 570203 540502
rect 583520 537692 584960 537932
rect 67633 537026 67699 537029
rect 67633 537024 70012 537026
rect 67633 536968 67638 537024
rect 67694 536968 70012 537024
rect 67633 536966 70012 536968
rect 67633 536963 67699 536966
rect 571701 532674 571767 532677
rect 569940 532672 571767 532674
rect 569940 532616 571706 532672
rect 571762 532616 571767 532672
rect 569940 532614 571767 532616
rect 571701 532611 571767 532614
rect 67449 529138 67515 529141
rect 67449 529136 70012 529138
rect 67449 529080 67454 529136
rect 67510 529080 70012 529136
rect 67449 529078 70012 529080
rect 67449 529075 67515 529078
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 571977 524786 572043 524789
rect 569940 524784 572043 524786
rect 569940 524728 571982 524784
rect 572038 524728 572043 524784
rect 569940 524726 572043 524728
rect 571977 524723 572043 524726
rect 580257 524514 580323 524517
rect 583520 524514 584960 524604
rect 580257 524512 584960 524514
rect 580257 524456 580262 524512
rect 580318 524456 584960 524512
rect 580257 524454 584960 524456
rect 580257 524451 580323 524454
rect 583520 524364 584960 524454
rect 67357 521250 67423 521253
rect 67357 521248 70012 521250
rect 67357 521192 67362 521248
rect 67418 521192 70012 521248
rect 67357 521190 70012 521192
rect 67357 521187 67423 521190
rect 570321 517170 570387 517173
rect 569940 517168 570387 517170
rect 569940 517112 570326 517168
rect 570382 517112 570387 517168
rect 569940 517110 570387 517112
rect 570321 517107 570387 517110
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 68737 513634 68803 513637
rect 68737 513632 70012 513634
rect 68737 513576 68742 513632
rect 68798 513576 70012 513632
rect 68737 513574 70012 513576
rect 68737 513571 68803 513574
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 572437 509282 572503 509285
rect 569940 509280 572503 509282
rect 569940 509224 572442 509280
rect 572498 509224 572503 509280
rect 569940 509222 572503 509224
rect 572437 509219 572503 509222
rect 67265 505746 67331 505749
rect 67265 505744 70012 505746
rect 67265 505688 67270 505744
rect 67326 505688 70012 505744
rect 67265 505686 70012 505688
rect 67265 505683 67331 505686
rect -960 501652 480 501892
rect 569358 500853 569418 501364
rect 569358 500848 569467 500853
rect 569358 500792 569406 500848
rect 569462 500792 569467 500848
rect 569358 500790 569467 500792
rect 569401 500787 569467 500790
rect 68645 497858 68711 497861
rect 68645 497856 70012 497858
rect 68645 497800 68650 497856
rect 68706 497800 70012 497856
rect 583520 497844 584960 498084
rect 68645 497798 70012 497800
rect 68645 497795 68711 497798
rect 569401 494050 569467 494053
rect 569358 494048 569467 494050
rect 569358 493992 569406 494048
rect 569462 493992 569467 494048
rect 569358 493987 569467 493992
rect 569358 493476 569418 493987
rect -960 488596 480 488836
rect 571425 485890 571491 485893
rect 569940 485888 571491 485890
rect 569940 485832 571430 485888
rect 571486 485832 571491 485888
rect 569940 485830 571491 485832
rect 571425 485827 571491 485830
rect 583520 484516 584960 484756
rect 68369 482354 68435 482357
rect 68369 482352 70012 482354
rect 68369 482296 68374 482352
rect 68430 482296 70012 482352
rect 68369 482294 70012 482296
rect 68369 482291 68435 482294
rect 571333 478002 571399 478005
rect 569940 478000 571399 478002
rect 569940 477944 571338 478000
rect 571394 477944 571399 478000
rect 569940 477942 571399 477944
rect 571333 477939 571399 477942
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 68277 474466 68343 474469
rect 68277 474464 70012 474466
rect 68277 474408 68282 474464
rect 68338 474408 70012 474464
rect 68277 474406 70012 474408
rect 68277 474403 68343 474406
rect 580257 471474 580323 471477
rect 583520 471474 584960 471564
rect 580257 471472 584960 471474
rect 580257 471416 580262 471472
rect 580318 471416 584960 471472
rect 580257 471414 584960 471416
rect 580257 471411 580323 471414
rect 583520 471324 584960 471414
rect 571517 470114 571583 470117
rect 569940 470112 571583 470114
rect 569940 470056 571522 470112
rect 571578 470056 571583 470112
rect 569940 470054 571583 470056
rect 571517 470051 571583 470054
rect 68553 466578 68619 466581
rect 68553 466576 70012 466578
rect 68553 466520 68558 466576
rect 68614 466520 70012 466576
rect 68553 466518 70012 466520
rect 68553 466515 68619 466518
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 570321 462498 570387 462501
rect 569940 462496 570387 462498
rect 569940 462440 570326 462496
rect 570382 462440 570387 462496
rect 569940 462438 570387 462440
rect 570321 462435 570387 462438
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 572621 454610 572687 454613
rect 569940 454608 572687 454610
rect 569940 454552 572626 454608
rect 572682 454552 572687 454608
rect 569940 454550 572687 454552
rect 572621 454547 572687 454550
rect 68645 451074 68711 451077
rect 68645 451072 70012 451074
rect 68645 451016 68650 451072
rect 68706 451016 70012 451072
rect 68645 451014 70012 451016
rect 68645 451011 68711 451014
rect -960 449428 480 449668
rect 569358 446181 569418 446692
rect 569358 446176 569467 446181
rect 569358 446120 569406 446176
rect 569462 446120 569467 446176
rect 569358 446118 569467 446120
rect 569401 446115 569467 446118
rect 583520 444668 584960 444908
rect 68461 443186 68527 443189
rect 68461 443184 70012 443186
rect 68461 443128 68466 443184
rect 68522 443128 70012 443184
rect 68461 443126 70012 443128
rect 68461 443123 68527 443126
rect -960 436508 480 436748
rect 67173 435298 67239 435301
rect 67173 435296 70012 435298
rect 67173 435240 67178 435296
rect 67234 435240 70012 435296
rect 67173 435238 70012 435240
rect 67173 435235 67239 435238
rect 569401 431490 569467 431493
rect 569358 431488 569467 431490
rect 569358 431432 569406 431488
rect 569462 431432 569467 431488
rect 583520 431476 584960 431716
rect 569358 431427 569467 431432
rect 569358 431188 569418 431427
rect 67909 427410 67975 427413
rect 67909 427408 70012 427410
rect 67909 427352 67914 427408
rect 67970 427352 70012 427408
rect 67909 427350 70012 427352
rect 67909 427347 67975 427350
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 570413 423330 570479 423333
rect 569940 423328 570479 423330
rect 569940 423272 570418 423328
rect 570474 423272 570479 423328
rect 569940 423270 570479 423272
rect 570413 423267 570479 423270
rect 67081 419794 67147 419797
rect 67081 419792 70012 419794
rect 67081 419736 67086 419792
rect 67142 419736 70012 419792
rect 67081 419734 70012 419736
rect 67081 419731 67147 419734
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 571609 415442 571675 415445
rect 569940 415440 571675 415442
rect 569940 415384 571614 415440
rect 571670 415384 571675 415440
rect 569940 415382 571675 415384
rect 571609 415379 571675 415382
rect 67633 411906 67699 411909
rect 67633 411904 70012 411906
rect 67633 411848 67638 411904
rect 67694 411848 70012 411904
rect 67633 411846 70012 411848
rect 67633 411843 67699 411846
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 570413 407554 570479 407557
rect 569940 407552 570479 407554
rect 569940 407496 570418 407552
rect 570474 407496 570479 407552
rect 569940 407494 570479 407496
rect 570413 407491 570479 407494
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 68001 404018 68067 404021
rect 68001 404016 70012 404018
rect 68001 403960 68006 404016
rect 68062 403960 70012 404016
rect 68001 403958 70012 403960
rect 68001 403955 68067 403958
rect 570505 399938 570571 399941
rect 569940 399936 570571 399938
rect 569940 399880 570510 399936
rect 570566 399880 570571 399936
rect 569940 399878 570571 399880
rect 570505 399875 570571 399878
rect -960 397340 480 397580
rect 67633 396402 67699 396405
rect 67633 396400 70012 396402
rect 67633 396344 67638 396400
rect 67694 396344 70012 396400
rect 67633 396342 70012 396344
rect 67633 396339 67699 396342
rect 572529 392050 572595 392053
rect 569940 392048 572595 392050
rect 569940 391992 572534 392048
rect 572590 391992 572595 392048
rect 569940 391990 572595 391992
rect 572529 391987 572595 391990
rect 583520 391628 584960 391868
rect 69013 388514 69079 388517
rect 69013 388512 70012 388514
rect 69013 388456 69018 388512
rect 69074 388456 70012 388512
rect 69013 388454 70012 388456
rect 69013 388451 69079 388454
rect -960 384284 480 384524
rect 571793 384162 571859 384165
rect 569940 384160 571859 384162
rect 569940 384104 571798 384160
rect 571854 384104 571859 384160
rect 569940 384102 571859 384104
rect 571793 384099 571859 384102
rect 583520 378300 584960 378540
rect 67633 372738 67699 372741
rect 67633 372736 70012 372738
rect 67633 372680 67638 372736
rect 67694 372680 70012 372736
rect 67633 372678 70012 372680
rect 67633 372675 67699 372678
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 67633 365122 67699 365125
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 67633 365120 70012 365122
rect 67633 365064 67638 365120
rect 67694 365064 70012 365120
rect 67633 365062 70012 365064
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 67633 365059 67699 365062
rect 579981 365059 580047 365062
rect 583520 364972 584960 365062
rect 572805 360770 572871 360773
rect 569940 360768 572871 360770
rect 569940 360712 572810 360768
rect 572866 360712 572871 360768
rect 569940 360710 572871 360712
rect 572805 360707 572871 360710
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 67817 357234 67883 357237
rect 67817 357232 70012 357234
rect 67817 357176 67822 357232
rect 67878 357176 70012 357232
rect 67817 357174 70012 357176
rect 67817 357171 67883 357174
rect 572897 352882 572963 352885
rect 569940 352880 572963 352882
rect 569940 352824 572902 352880
rect 572958 352824 572963 352880
rect 569940 352822 572963 352824
rect 572897 352819 572963 352822
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 67633 349346 67699 349349
rect 67633 349344 70012 349346
rect 67633 349288 67638 349344
rect 67694 349288 70012 349344
rect 67633 349286 70012 349288
rect 67633 349283 67699 349286
rect -960 345252 480 345492
rect 572069 344994 572135 344997
rect 569940 344992 572135 344994
rect 569940 344936 572074 344992
rect 572130 344936 572135 344992
rect 569940 344934 572135 344936
rect 572069 344931 572135 344934
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 572621 329490 572687 329493
rect 569940 329488 572687 329490
rect 569940 329432 572626 329488
rect 572682 329432 572687 329488
rect 569940 329430 572687 329432
rect 572621 329427 572687 329430
rect 67633 325954 67699 325957
rect 67633 325952 70012 325954
rect 67633 325896 67638 325952
rect 67694 325896 70012 325952
rect 67633 325894 70012 325896
rect 67633 325891 67699 325894
rect 583520 325124 584960 325364
rect 569309 321874 569375 321877
rect 569309 321872 569418 321874
rect 569309 321816 569314 321872
rect 569370 321816 569418 321872
rect 569309 321811 569418 321816
rect 569358 321572 569418 321811
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 69197 318066 69263 318069
rect 69197 318064 70012 318066
rect 69197 318008 69202 318064
rect 69258 318008 70012 318064
rect 69197 318006 70012 318008
rect 69197 318003 69263 318006
rect 580349 312082 580415 312085
rect 583520 312082 584960 312172
rect 580349 312080 584960 312082
rect 580349 312024 580354 312080
rect 580410 312024 584960 312080
rect 580349 312022 584960 312024
rect 580349 312019 580415 312022
rect 583520 311932 584960 312022
rect 69105 310178 69171 310181
rect 69105 310176 70012 310178
rect 69105 310120 69110 310176
rect 69166 310120 70012 310176
rect 69105 310118 70012 310120
rect 69105 310115 69171 310118
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 571333 306098 571399 306101
rect 569940 306096 571399 306098
rect 569940 306040 571338 306096
rect 571394 306040 571399 306096
rect 569940 306038 571399 306040
rect 571333 306035 571399 306038
rect 67817 302562 67883 302565
rect 67817 302560 70012 302562
rect 67817 302504 67822 302560
rect 67878 302504 70012 302560
rect 67817 302502 70012 302504
rect 67817 302499 67883 302502
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 571885 298210 571951 298213
rect 569940 298208 571951 298210
rect 569940 298152 571890 298208
rect 571946 298152 571951 298208
rect 569940 298150 571951 298152
rect 571885 298147 571951 298150
rect 69289 294674 69355 294677
rect 69289 294672 70012 294674
rect 69289 294616 69294 294672
rect 69350 294616 70012 294672
rect 69289 294614 70012 294616
rect 69289 294611 69355 294614
rect -960 293028 480 293268
rect 67817 286786 67883 286789
rect 67817 286784 70012 286786
rect 67817 286728 67822 286784
rect 67878 286728 70012 286784
rect 67817 286726 70012 286728
rect 67817 286723 67883 286726
rect 583520 285276 584960 285516
rect 571977 282706 572043 282709
rect 569940 282704 572043 282706
rect 569940 282648 571982 282704
rect 572038 282648 572043 282704
rect 569940 282646 572043 282648
rect 571977 282643 572043 282646
rect -960 279972 480 280212
rect 68185 278898 68251 278901
rect 68185 278896 70012 278898
rect 68185 278840 68190 278896
rect 68246 278840 70012 278896
rect 68185 278838 70012 278840
rect 68185 278835 68251 278838
rect 570597 274818 570663 274821
rect 569940 274816 570663 274818
rect 569940 274760 570602 274816
rect 570658 274760 570663 274816
rect 569940 274758 570663 274760
rect 570597 274755 570663 274758
rect 583520 272084 584960 272324
rect 67633 271282 67699 271285
rect 67633 271280 70012 271282
rect 67633 271224 67638 271280
rect 67694 271224 70012 271280
rect 67633 271222 70012 271224
rect 67633 271219 67699 271222
rect -960 267202 480 267292
rect 3785 267202 3851 267205
rect -960 267200 3851 267202
rect -960 267144 3790 267200
rect 3846 267144 3851 267200
rect -960 267142 3851 267144
rect -960 267052 480 267142
rect 3785 267139 3851 267142
rect 569358 266525 569418 266900
rect 569309 266520 569418 266525
rect 569309 266464 569314 266520
rect 569370 266464 569418 266520
rect 569309 266462 569418 266464
rect 569309 266459 569375 266462
rect 68277 263394 68343 263397
rect 68277 263392 70012 263394
rect 68277 263336 68282 263392
rect 68338 263336 70012 263392
rect 68277 263334 70012 263336
rect 68277 263331 68343 263334
rect 569358 258637 569418 259012
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect 569309 258632 569418 258637
rect 569309 258576 569314 258632
rect 569370 258576 569418 258632
rect 569309 258574 569418 258576
rect 569309 258571 569375 258574
rect 68185 255506 68251 255509
rect 68185 255504 70012 255506
rect 68185 255448 68190 255504
rect 68246 255448 70012 255504
rect 68185 255446 70012 255448
rect 68185 255443 68251 255446
rect -960 254146 480 254236
rect 4061 254146 4127 254149
rect -960 254144 4127 254146
rect -960 254088 4066 254144
rect 4122 254088 4127 254144
rect -960 254086 4127 254088
rect -960 253996 480 254086
rect 4061 254083 4127 254086
rect 572069 251426 572135 251429
rect 569940 251424 572135 251426
rect 569940 251368 572074 251424
rect 572130 251368 572135 251424
rect 569940 251366 572135 251368
rect 572069 251363 572135 251366
rect 68369 247618 68435 247621
rect 68369 247616 70012 247618
rect 68369 247560 68374 247616
rect 68430 247560 70012 247616
rect 68369 247558 70012 247560
rect 68369 247555 68435 247558
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 569542 242861 569602 243508
rect 569542 242856 569651 242861
rect 569542 242800 569590 242856
rect 569646 242800 569651 242856
rect 569542 242798 569651 242800
rect 569585 242795 569651 242798
rect -960 240940 480 241180
rect 67633 240002 67699 240005
rect 67633 240000 70012 240002
rect 67633 239944 67638 240000
rect 67694 239944 70012 240000
rect 67633 239942 70012 239944
rect 67633 239939 67699 239942
rect 569358 235109 569418 235620
rect 569309 235104 569418 235109
rect 569309 235048 569314 235104
rect 569370 235048 569418 235104
rect 569309 235046 569418 235048
rect 569309 235043 569375 235046
rect 583520 232236 584960 232476
rect 67633 232114 67699 232117
rect 67633 232112 70012 232114
rect 67633 232056 67638 232112
rect 67694 232056 70012 232112
rect 67633 232054 70012 232056
rect 67633 232051 67699 232054
rect -960 227884 480 228124
rect 572161 227762 572227 227765
rect 569940 227760 572227 227762
rect 569940 227704 572166 227760
rect 572222 227704 572227 227760
rect 569940 227702 572227 227704
rect 572161 227699 572227 227702
rect 66989 224226 67055 224229
rect 66989 224224 70012 224226
rect 66989 224168 66994 224224
rect 67050 224168 70012 224224
rect 66989 224166 70012 224168
rect 66989 224163 67055 224166
rect 569358 219877 569418 220116
rect 569358 219872 569467 219877
rect 569358 219816 569406 219872
rect 569462 219816 569467 219872
rect 569358 219814 569467 219816
rect 569401 219811 569467 219814
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3233 214978 3299 214981
rect -960 214976 3299 214978
rect -960 214920 3238 214976
rect 3294 214920 3299 214976
rect -960 214918 3299 214920
rect -960 214828 480 214918
rect 3233 214915 3299 214918
rect 570689 212258 570755 212261
rect 569940 212256 570755 212258
rect 569940 212200 570694 212256
rect 570750 212200 570755 212256
rect 569940 212198 570755 212200
rect 570689 212195 570755 212198
rect 67633 208722 67699 208725
rect 67633 208720 70012 208722
rect 67633 208664 67638 208720
rect 67694 208664 70012 208720
rect 67633 208662 70012 208664
rect 67633 208659 67699 208662
rect 580441 205730 580507 205733
rect 583520 205730 584960 205820
rect 580441 205728 584960 205730
rect 580441 205672 580446 205728
rect 580502 205672 584960 205728
rect 580441 205670 584960 205672
rect 580441 205667 580507 205670
rect 583520 205580 584960 205670
rect 569358 204101 569418 204340
rect 569358 204096 569467 204101
rect 569358 204040 569406 204096
rect 569462 204040 569467 204096
rect 569358 204038 569467 204040
rect 569401 204035 569467 204038
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 67725 200834 67791 200837
rect 67725 200832 70012 200834
rect 67725 200776 67730 200832
rect 67786 200776 70012 200832
rect 67725 200774 70012 200776
rect 67725 200771 67791 200774
rect 570873 196482 570939 196485
rect 569940 196480 570939 196482
rect 569940 196424 570878 196480
rect 570934 196424 570939 196480
rect 569940 196422 570939 196424
rect 570873 196419 570939 196422
rect 68093 192946 68159 192949
rect 68093 192944 70012 192946
rect 68093 192888 68098 192944
rect 68154 192888 70012 192944
rect 68093 192886 70012 192888
rect 68093 192883 68159 192886
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 570965 188866 571031 188869
rect 569940 188864 571031 188866
rect 569940 188808 570970 188864
rect 571026 188808 571031 188864
rect 569940 188806 571031 188808
rect 570965 188803 571031 188806
rect 66897 185330 66963 185333
rect 66897 185328 70012 185330
rect 66897 185272 66902 185328
rect 66958 185272 70012 185328
rect 66897 185270 70012 185272
rect 66897 185267 66963 185270
rect 579889 179210 579955 179213
rect 583520 179210 584960 179300
rect 579889 179208 584960 179210
rect 579889 179152 579894 179208
rect 579950 179152 584960 179208
rect 579889 179150 584960 179152
rect 579889 179147 579955 179150
rect 583520 179060 584960 179150
rect 67633 177442 67699 177445
rect 67633 177440 70012 177442
rect 67633 177384 67638 177440
rect 67694 177384 70012 177440
rect 67633 177382 70012 177384
rect 67633 177379 67699 177382
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 570229 165202 570295 165205
rect 569940 165200 570295 165202
rect 569940 165144 570234 165200
rect 570290 165144 570295 165200
rect 569940 165142 570295 165144
rect 570229 165139 570295 165142
rect -960 162890 480 162980
rect 3693 162890 3759 162893
rect -960 162888 3759 162890
rect -960 162832 3698 162888
rect 3754 162832 3759 162888
rect -960 162830 3759 162832
rect -960 162740 480 162830
rect 3693 162827 3759 162830
rect 67633 161666 67699 161669
rect 67633 161664 70012 161666
rect 67633 161608 67638 161664
rect 67694 161608 70012 161664
rect 67633 161606 70012 161608
rect 67633 161603 67699 161606
rect 570045 158130 570111 158133
rect 569910 158128 570111 158130
rect 569910 158072 570050 158128
rect 570106 158072 570111 158128
rect 569910 158070 570111 158072
rect 569910 157556 569970 158070
rect 570045 158067 570111 158070
rect 68001 154050 68067 154053
rect 68001 154048 70012 154050
rect 68001 153992 68006 154048
rect 68062 153992 70012 154048
rect 68001 153990 70012 153992
rect 68001 153987 68067 153990
rect 583520 152540 584960 152780
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 569542 149157 569602 149668
rect 569493 149152 569602 149157
rect 569493 149096 569498 149152
rect 569554 149096 569602 149152
rect 569493 149094 569602 149096
rect 569493 149091 569559 149094
rect 67909 146162 67975 146165
rect 67909 146160 70012 146162
rect 67909 146104 67914 146160
rect 67970 146104 70012 146160
rect 67909 146102 70012 146104
rect 67909 146099 67975 146102
rect 571701 141810 571767 141813
rect 569940 141808 571767 141810
rect 569940 141752 571706 141808
rect 571762 141752 571767 141808
rect 569940 141750 571767 141752
rect 571701 141747 571767 141750
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 67633 138274 67699 138277
rect 67633 138272 70012 138274
rect 67633 138216 67638 138272
rect 67694 138216 70012 138272
rect 67633 138214 70012 138216
rect 67633 138211 67699 138214
rect -960 136628 480 136868
rect 569910 133922 569970 134164
rect 570045 133922 570111 133925
rect 569910 133920 570111 133922
rect 569910 133864 570050 133920
rect 570106 133864 570111 133920
rect 569910 133862 570111 133864
rect 570045 133859 570111 133862
rect 67633 130386 67699 130389
rect 67633 130384 70012 130386
rect 67633 130328 67638 130384
rect 67694 130328 70012 130384
rect 67633 130326 70012 130328
rect 67633 130323 67699 130326
rect 569953 126850 570019 126853
rect 569910 126848 570019 126850
rect 569910 126792 569958 126848
rect 570014 126792 570019 126848
rect 569910 126787 570019 126792
rect 569910 126276 569970 126787
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 68093 122770 68159 122773
rect 68093 122768 70012 122770
rect 68093 122712 68098 122768
rect 68154 122712 70012 122768
rect 68093 122710 70012 122712
rect 68093 122707 68159 122710
rect 569726 117877 569786 118388
rect 569677 117872 569786 117877
rect 569677 117816 569682 117872
rect 569738 117816 569786 117872
rect 569677 117814 569786 117816
rect 569677 117811 569743 117814
rect 67817 114882 67883 114885
rect 67817 114880 70012 114882
rect 67817 114824 67822 114880
rect 67878 114824 70012 114880
rect 67817 114822 70012 114824
rect 67817 114819 67883 114822
rect 583520 112692 584960 112932
rect -960 110666 480 110756
rect 3601 110666 3667 110669
rect -960 110664 3667 110666
rect -960 110608 3606 110664
rect 3662 110608 3667 110664
rect -960 110606 3667 110608
rect -960 110516 480 110606
rect 3601 110603 3667 110606
rect 572253 110530 572319 110533
rect 569940 110528 572319 110530
rect 569940 110472 572258 110528
rect 572314 110472 572319 110528
rect 569940 110470 572319 110472
rect 572253 110467 572319 110470
rect 572345 102914 572411 102917
rect 569940 102912 572411 102914
rect 569940 102856 572350 102912
rect 572406 102856 572411 102912
rect 569940 102854 572411 102856
rect 572345 102851 572411 102854
rect 579705 99514 579771 99517
rect 583520 99514 584960 99604
rect 579705 99512 584960 99514
rect 579705 99456 579710 99512
rect 579766 99456 584960 99512
rect 579705 99454 584960 99456
rect 579705 99451 579771 99454
rect 583520 99364 584960 99454
rect 67633 99106 67699 99109
rect 67633 99104 70012 99106
rect 67633 99048 67638 99104
rect 67694 99048 70012 99104
rect 67633 99046 70012 99048
rect 67633 99043 67699 99046
rect -960 97610 480 97700
rect 3325 97610 3391 97613
rect -960 97608 3391 97610
rect -960 97552 3330 97608
rect 3386 97552 3391 97608
rect -960 97550 3391 97552
rect -960 97460 480 97550
rect 3325 97547 3391 97550
rect 570229 95026 570295 95029
rect 569940 95024 570295 95026
rect 569940 94968 570234 95024
rect 570290 94968 570295 95024
rect 569940 94966 570295 94968
rect 570229 94963 570295 94966
rect 67633 91490 67699 91493
rect 67633 91488 70012 91490
rect 67633 91432 67638 91488
rect 67694 91432 70012 91488
rect 67633 91430 70012 91432
rect 67633 91427 67699 91430
rect 569953 87410 570019 87413
rect 569910 87408 570019 87410
rect 569910 87352 569958 87408
rect 570014 87352 570019 87408
rect 569910 87347 570019 87352
rect 569910 87108 569970 87347
rect 580533 86186 580599 86189
rect 583520 86186 584960 86276
rect 580533 86184 584960 86186
rect 580533 86128 580538 86184
rect 580594 86128 584960 86184
rect 580533 86126 584960 86128
rect 580533 86123 580599 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 68369 83602 68435 83605
rect 68369 83600 70012 83602
rect 68369 83544 68374 83600
rect 68430 83544 70012 83600
rect 68369 83542 70012 83544
rect 68369 83539 68435 83542
rect 571333 79250 571399 79253
rect 569940 79248 571399 79250
rect 569940 79192 571338 79248
rect 571394 79192 571399 79248
rect 569940 79190 571399 79192
rect 571333 79187 571399 79190
rect 583520 72844 584960 73084
rect -960 71634 480 71724
rect 3877 71634 3943 71637
rect -960 71632 3943 71634
rect -960 71576 3882 71632
rect 3938 71576 3943 71632
rect -960 71574 3943 71576
rect -960 71484 480 71574
rect 3877 71571 3943 71574
rect 569358 71093 569418 71604
rect 569309 71088 569418 71093
rect 569309 71032 569314 71088
rect 569370 71032 569418 71088
rect 569309 71030 569418 71032
rect 569309 71027 569375 71030
rect 223297 67554 223363 67557
rect 429142 67554 429148 67556
rect 223297 67552 429148 67554
rect 223297 67496 223302 67552
rect 223358 67496 429148 67552
rect 223297 67494 429148 67496
rect 223297 67491 223363 67494
rect 429142 67492 429148 67494
rect 429212 67492 429218 67556
rect 106774 67356 106780 67420
rect 106844 67418 106850 67420
rect 307937 67418 308003 67421
rect 106844 67416 308003 67418
rect 106844 67360 307942 67416
rect 307998 67360 308003 67416
rect 106844 67358 308003 67360
rect 106844 67356 106850 67358
rect 307937 67355 308003 67358
rect 180977 67282 181043 67285
rect 234654 67282 234660 67284
rect 180977 67280 234660 67282
rect 180977 67224 180982 67280
rect 181038 67224 234660 67280
rect 180977 67222 234660 67224
rect 180977 67219 181043 67222
rect 234654 67220 234660 67222
rect 234724 67220 234730 67284
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580349 46338 580415 46341
rect 583520 46338 584960 46428
rect 580349 46336 584960 46338
rect 580349 46280 580354 46336
rect 580410 46280 584960 46336
rect 580349 46278 584960 46280
rect 580349 46275 580415 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32466 480 32556
rect 3693 32466 3759 32469
rect -960 32464 3759 32466
rect -960 32408 3698 32464
rect 3754 32408 3759 32464
rect -960 32406 3759 32408
rect -960 32316 480 32406
rect 3693 32403 3759 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 226333 6898 226399 6901
rect 346894 6898 346900 6900
rect 226333 6896 346900 6898
rect 226333 6840 226338 6896
rect 226394 6840 346900 6896
rect 226333 6838 346900 6840
rect 226333 6835 226399 6838
rect 346894 6836 346900 6838
rect 346964 6836 346970 6900
rect 150617 6762 150683 6765
rect 345054 6762 345060 6764
rect 150617 6760 345060 6762
rect 150617 6704 150622 6760
rect 150678 6704 345060 6760
rect 150617 6702 345060 6704
rect 150617 6699 150683 6702
rect 345054 6700 345060 6702
rect 345124 6700 345130 6764
rect 200297 6626 200363 6629
rect 403566 6626 403572 6628
rect 200297 6624 403572 6626
rect -960 6340 480 6580
rect 200297 6568 200302 6624
rect 200358 6568 403572 6624
rect 200297 6566 403572 6568
rect 200297 6563 200363 6566
rect 403566 6564 403572 6566
rect 403636 6564 403642 6628
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 101990 6428 101996 6492
rect 102060 6490 102066 6492
rect 233417 6490 233483 6493
rect 102060 6488 233483 6490
rect 102060 6432 233422 6488
rect 233478 6432 233483 6488
rect 102060 6430 233483 6432
rect 102060 6428 102066 6430
rect 233417 6427 233483 6430
rect 237005 6490 237071 6493
rect 460974 6490 460980 6492
rect 237005 6488 460980 6490
rect 237005 6432 237010 6488
rect 237066 6432 460980 6488
rect 237005 6430 460980 6432
rect 237005 6427 237071 6430
rect 460974 6428 460980 6430
rect 461044 6428 461050 6492
rect 583520 6476 584960 6566
rect 195605 6354 195671 6357
rect 440182 6354 440188 6356
rect 195605 6352 440188 6354
rect 195605 6296 195610 6352
rect 195666 6296 440188 6352
rect 195605 6294 440188 6296
rect 195605 6291 195671 6294
rect 440182 6292 440188 6294
rect 440252 6292 440258 6356
rect 180241 6218 180307 6221
rect 481766 6218 481772 6220
rect 180241 6216 481772 6218
rect 180241 6160 180246 6216
rect 180302 6160 481772 6216
rect 180241 6158 481772 6160
rect 180241 6155 180307 6158
rect 481766 6156 481772 6158
rect 481836 6156 481842 6220
rect 183737 6082 183803 6085
rect 281574 6082 281580 6084
rect 183737 6080 281580 6082
rect 183737 6024 183742 6080
rect 183798 6024 281580 6080
rect 183737 6022 281580 6024
rect 183737 6019 183803 6022
rect 281574 6020 281580 6022
rect 281644 6020 281650 6084
rect 161289 5946 161355 5949
rect 244222 5946 244228 5948
rect 161289 5944 244228 5946
rect 161289 5888 161294 5944
rect 161350 5888 244228 5944
rect 161289 5886 244228 5888
rect 161289 5883 161355 5886
rect 244222 5884 244228 5886
rect 244292 5884 244298 5948
rect 133638 5476 133644 5540
rect 133708 5538 133714 5540
rect 166073 5538 166139 5541
rect 133708 5536 166139 5538
rect 133708 5480 166078 5536
rect 166134 5480 166139 5536
rect 133708 5478 166139 5480
rect 133708 5476 133714 5478
rect 166073 5475 166139 5478
rect 144678 5340 144684 5404
rect 144748 5402 144754 5404
rect 201493 5402 201559 5405
rect 144748 5400 201559 5402
rect 144748 5344 201498 5400
rect 201554 5344 201559 5400
rect 144748 5342 201559 5344
rect 144748 5340 144754 5342
rect 201493 5339 201559 5342
rect 109309 5266 109375 5269
rect 175774 5266 175780 5268
rect 109309 5264 175780 5266
rect 109309 5208 109314 5264
rect 109370 5208 175780 5264
rect 109309 5206 175780 5208
rect 109309 5203 109375 5206
rect 175774 5204 175780 5206
rect 175844 5204 175850 5268
rect 203885 5266 203951 5269
rect 270534 5266 270540 5268
rect 203885 5264 270540 5266
rect 203885 5208 203890 5264
rect 203946 5208 270540 5264
rect 203885 5206 270540 5208
rect 203885 5203 203951 5206
rect 270534 5204 270540 5206
rect 270604 5204 270610 5268
rect 86718 5068 86724 5132
rect 86788 5130 86794 5132
rect 135253 5130 135319 5133
rect 86788 5128 135319 5130
rect 86788 5072 135258 5128
rect 135314 5072 135319 5128
rect 86788 5070 135319 5072
rect 86788 5068 86794 5070
rect 135253 5067 135319 5070
rect 155718 5068 155724 5132
rect 155788 5130 155794 5132
rect 168373 5130 168439 5133
rect 155788 5128 168439 5130
rect 155788 5072 168378 5128
rect 168434 5072 168439 5128
rect 155788 5070 168439 5072
rect 155788 5068 155794 5070
rect 168373 5067 168439 5070
rect 170990 5068 170996 5132
rect 171060 5130 171066 5132
rect 238109 5130 238175 5133
rect 171060 5128 238175 5130
rect 171060 5072 238114 5128
rect 238170 5072 238175 5128
rect 171060 5070 238175 5072
rect 171060 5068 171066 5070
rect 238109 5067 238175 5070
rect 108113 4994 108179 4997
rect 168966 4994 168972 4996
rect 108113 4992 168972 4994
rect 108113 4936 108118 4992
rect 108174 4936 168972 4992
rect 108113 4934 168972 4936
rect 108113 4931 108179 4934
rect 168966 4932 168972 4934
rect 169036 4932 169042 4996
rect 170765 4994 170831 4997
rect 348366 4994 348372 4996
rect 170765 4992 348372 4994
rect 170765 4936 170770 4992
rect 170826 4936 348372 4992
rect 170765 4934 348372 4936
rect 170765 4931 170831 4934
rect 348366 4932 348372 4934
rect 348436 4932 348442 4996
rect 118785 4858 118851 4861
rect 550766 4858 550772 4860
rect 118785 4856 550772 4858
rect 118785 4800 118790 4856
rect 118846 4800 550772 4856
rect 118785 4798 550772 4800
rect 118785 4795 118851 4798
rect 550766 4796 550772 4798
rect 550836 4796 550842 4860
rect 130561 3770 130627 3773
rect 130878 3770 130884 3772
rect 130561 3768 130884 3770
rect 130561 3712 130566 3768
rect 130622 3712 130884 3768
rect 130561 3710 130884 3712
rect 130561 3707 130627 3710
rect 130878 3708 130884 3710
rect 130948 3708 130954 3772
rect 140037 3770 140103 3773
rect 140630 3770 140636 3772
rect 140037 3768 140636 3770
rect 140037 3712 140042 3768
rect 140098 3712 140636 3768
rect 140037 3710 140636 3712
rect 140037 3707 140103 3710
rect 140630 3708 140636 3710
rect 140700 3708 140706 3772
rect 145598 3708 145604 3772
rect 145668 3770 145674 3772
rect 145925 3770 145991 3773
rect 153009 3772 153075 3773
rect 145668 3768 145991 3770
rect 145668 3712 145930 3768
rect 145986 3712 145991 3768
rect 145668 3710 145991 3712
rect 145668 3708 145674 3710
rect 145925 3707 145991 3710
rect 152958 3708 152964 3772
rect 153028 3770 153075 3772
rect 156597 3772 156663 3773
rect 156597 3770 156644 3772
rect 153028 3768 153120 3770
rect 153070 3712 153120 3768
rect 153028 3710 153120 3712
rect 156552 3768 156644 3770
rect 156552 3712 156602 3768
rect 156552 3710 156644 3712
rect 153028 3708 153075 3710
rect 153009 3707 153075 3708
rect 156597 3708 156644 3710
rect 156708 3708 156714 3772
rect 160093 3770 160159 3773
rect 161238 3770 161244 3772
rect 160093 3768 161244 3770
rect 160093 3712 160098 3768
rect 160154 3712 161244 3768
rect 160093 3710 161244 3712
rect 156597 3707 156663 3708
rect 160093 3707 160159 3710
rect 161238 3708 161244 3710
rect 161308 3708 161314 3772
rect 164550 3708 164556 3772
rect 164620 3770 164626 3772
rect 164877 3770 164943 3773
rect 164620 3768 164943 3770
rect 164620 3712 164882 3768
rect 164938 3712 164943 3768
rect 164620 3710 164943 3712
rect 164620 3708 164626 3710
rect 164877 3707 164943 3710
rect 106917 3634 106983 3637
rect 117589 3634 117655 3637
rect 177982 3634 177988 3636
rect 106917 3632 113190 3634
rect 106917 3576 106922 3632
rect 106978 3576 113190 3632
rect 106917 3574 113190 3576
rect 106917 3571 106983 3574
rect 92749 3498 92815 3501
rect 93710 3498 93716 3500
rect 92749 3496 93716 3498
rect 92749 3440 92754 3496
rect 92810 3440 93716 3496
rect 92749 3438 93716 3440
rect 92749 3435 92815 3438
rect 93710 3436 93716 3438
rect 93780 3436 93786 3500
rect 97441 3498 97507 3501
rect 97758 3498 97764 3500
rect 97441 3496 97764 3498
rect 97441 3440 97446 3496
rect 97502 3440 97764 3496
rect 97441 3438 97764 3440
rect 97441 3435 97507 3438
rect 97758 3436 97764 3438
rect 97828 3436 97834 3500
rect 110505 3498 110571 3501
rect 111558 3498 111564 3500
rect 110505 3496 111564 3498
rect 110505 3440 110510 3496
rect 110566 3440 111564 3496
rect 110505 3438 111564 3440
rect 110505 3435 110571 3438
rect 111558 3436 111564 3438
rect 111628 3436 111634 3500
rect 113130 3498 113190 3574
rect 117589 3632 177988 3634
rect 117589 3576 117594 3632
rect 117650 3576 177988 3632
rect 117589 3574 177988 3576
rect 117589 3571 117655 3574
rect 177982 3572 177988 3574
rect 178052 3572 178058 3636
rect 205081 3634 205147 3637
rect 205398 3634 205404 3636
rect 205081 3632 205404 3634
rect 205081 3576 205086 3632
rect 205142 3576 205404 3632
rect 205081 3574 205404 3576
rect 205081 3571 205147 3574
rect 205398 3572 205404 3574
rect 205468 3572 205474 3636
rect 210969 3634 211035 3637
rect 214414 3634 214420 3636
rect 210969 3632 214420 3634
rect 210969 3576 210974 3632
rect 211030 3576 214420 3632
rect 210969 3574 214420 3576
rect 210969 3571 211035 3574
rect 214414 3572 214420 3574
rect 214484 3572 214490 3636
rect 220445 3634 220511 3637
rect 227529 3636 227595 3637
rect 220670 3634 220676 3636
rect 220445 3632 220676 3634
rect 220445 3576 220450 3632
rect 220506 3576 220676 3632
rect 220445 3574 220676 3576
rect 220445 3571 220511 3574
rect 220670 3572 220676 3574
rect 220740 3572 220746 3636
rect 227478 3572 227484 3636
rect 227548 3634 227595 3636
rect 227548 3632 227640 3634
rect 227590 3576 227640 3632
rect 227548 3574 227640 3576
rect 227548 3572 227595 3574
rect 227529 3571 227595 3572
rect 386454 3498 386460 3500
rect 113130 3438 386460 3498
rect 386454 3436 386460 3438
rect 386524 3436 386530 3500
rect 105721 3362 105787 3365
rect 539542 3362 539548 3364
rect 105721 3360 539548 3362
rect 105721 3304 105726 3360
rect 105782 3304 539548 3360
rect 105721 3302 539548 3304
rect 105721 3299 105787 3302
rect 539542 3300 539548 3302
rect 539612 3300 539618 3364
<< via3 >>
rect 106780 699756 106844 699820
rect 234660 699756 234724 699820
rect 429148 699756 429212 699820
rect 152964 571236 153028 571300
rect 175780 571100 175844 571164
rect 156644 570964 156708 571028
rect 227484 570964 227548 571028
rect 111564 570828 111628 570892
rect 346900 570828 346964 570892
rect 93716 570692 93780 570756
rect 348372 570692 348436 570756
rect 97764 570556 97828 570620
rect 168972 570420 169036 570484
rect 161244 570284 161308 570348
rect 145604 570148 145668 570212
rect 403572 570148 403636 570212
rect 220676 570012 220740 570076
rect 177988 568516 178052 568580
rect 86724 567292 86788 567356
rect 101996 567352 102060 567356
rect 101996 567296 102046 567352
rect 102046 567296 102060 567352
rect 101996 567292 102060 567296
rect 133644 567292 133708 567356
rect 144684 567292 144748 567356
rect 155724 567292 155788 567356
rect 170996 567352 171060 567356
rect 170996 567296 171010 567352
rect 171010 567296 171060 567352
rect 170996 567292 171060 567296
rect 210372 567292 210436 567356
rect 214420 567156 214484 567220
rect 244228 567292 244292 567356
rect 270540 567292 270604 567356
rect 281580 567292 281644 567356
rect 328500 567292 328564 567356
rect 345060 567292 345124 567356
rect 386460 567292 386524 567356
rect 440188 567292 440252 567356
rect 460980 567292 461044 567356
rect 481772 567292 481836 567356
rect 539548 567292 539612 567356
rect 550772 567292 550836 567356
rect 164556 566612 164620 566676
rect 130884 566476 130948 566540
rect 328500 566476 328564 566540
rect 140636 566340 140700 566404
rect 205404 565932 205468 565996
rect 210372 565932 210436 565996
rect 429148 67492 429212 67556
rect 106780 67356 106844 67420
rect 234660 67220 234724 67284
rect 346900 6836 346964 6900
rect 345060 6700 345124 6764
rect 403572 6564 403636 6628
rect 101996 6428 102060 6492
rect 460980 6428 461044 6492
rect 440188 6292 440252 6356
rect 481772 6156 481836 6220
rect 281580 6020 281644 6084
rect 244228 5884 244292 5948
rect 133644 5476 133708 5540
rect 144684 5340 144748 5404
rect 175780 5204 175844 5268
rect 270540 5204 270604 5268
rect 86724 5068 86788 5132
rect 155724 5068 155788 5132
rect 170996 5068 171060 5132
rect 168972 4932 169036 4996
rect 348372 4932 348436 4996
rect 550772 4796 550836 4860
rect 130884 3708 130948 3772
rect 140636 3708 140700 3772
rect 145604 3708 145668 3772
rect 152964 3768 153028 3772
rect 152964 3712 153014 3768
rect 153014 3712 153028 3768
rect 152964 3708 153028 3712
rect 156644 3768 156708 3772
rect 156644 3712 156658 3768
rect 156658 3712 156708 3768
rect 156644 3708 156708 3712
rect 161244 3708 161308 3772
rect 164556 3708 164620 3772
rect 93716 3436 93780 3500
rect 97764 3436 97828 3500
rect 111564 3436 111628 3500
rect 177988 3572 178052 3636
rect 205404 3572 205468 3636
rect 214420 3572 214484 3636
rect 220676 3572 220740 3636
rect 227484 3632 227548 3636
rect 227484 3576 227534 3632
rect 227534 3576 227548 3632
rect 227484 3572 227548 3576
rect 386460 3436 386524 3500
rect 539548 3300 539612 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 570000 74414 578898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 570000 78134 582618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 570000 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 570000 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 570000 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 93715 570756 93781 570757
rect 93715 570692 93716 570756
rect 93780 570692 93781 570756
rect 93715 570691 93781 570692
rect 86723 567356 86789 567357
rect 86723 567292 86724 567356
rect 86788 567292 86789 567356
rect 86723 567291 86789 567292
rect 74208 543454 74528 543486
rect 74208 543218 74250 543454
rect 74486 543218 74528 543454
rect 74208 543134 74528 543218
rect 74208 542898 74250 543134
rect 74486 542898 74528 543134
rect 74208 542866 74528 542898
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 74208 507454 74528 507486
rect 74208 507218 74250 507454
rect 74486 507218 74528 507454
rect 74208 507134 74528 507218
rect 74208 506898 74250 507134
rect 74486 506898 74528 507134
rect 74208 506866 74528 506898
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 74208 471454 74528 471486
rect 74208 471218 74250 471454
rect 74486 471218 74528 471454
rect 74208 471134 74528 471218
rect 74208 470898 74250 471134
rect 74486 470898 74528 471134
rect 74208 470866 74528 470898
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 74208 435454 74528 435486
rect 74208 435218 74250 435454
rect 74486 435218 74528 435454
rect 74208 435134 74528 435218
rect 74208 434898 74250 435134
rect 74486 434898 74528 435134
rect 74208 434866 74528 434898
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 74208 399454 74528 399486
rect 74208 399218 74250 399454
rect 74486 399218 74528 399454
rect 74208 399134 74528 399218
rect 74208 398898 74250 399134
rect 74486 398898 74528 399134
rect 74208 398866 74528 398898
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 74208 327454 74528 327486
rect 74208 327218 74250 327454
rect 74486 327218 74528 327454
rect 74208 327134 74528 327218
rect 74208 326898 74250 327134
rect 74486 326898 74528 327134
rect 74208 326866 74528 326898
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 74208 291454 74528 291486
rect 74208 291218 74250 291454
rect 74486 291218 74528 291454
rect 74208 291134 74528 291218
rect 74208 290898 74250 291134
rect 74486 290898 74528 291134
rect 74208 290866 74528 290898
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 74208 219454 74528 219486
rect 74208 219218 74250 219454
rect 74486 219218 74528 219454
rect 74208 219134 74528 219218
rect 74208 218898 74250 219134
rect 74486 218898 74528 219134
rect 74208 218866 74528 218898
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 74208 183454 74528 183486
rect 74208 183218 74250 183454
rect 74486 183218 74528 183454
rect 74208 183134 74528 183218
rect 74208 182898 74250 183134
rect 74486 182898 74528 183134
rect 74208 182866 74528 182898
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 74208 147454 74528 147486
rect 74208 147218 74250 147454
rect 74486 147218 74528 147454
rect 74208 147134 74528 147218
rect 74208 146898 74250 147134
rect 74486 146898 74528 147134
rect 74208 146866 74528 146898
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 74208 111454 74528 111486
rect 74208 111218 74250 111454
rect 74486 111218 74528 111454
rect 74208 111134 74528 111218
rect 74208 110898 74250 111134
rect 74486 110898 74528 111134
rect 74208 110866 74528 110898
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 74208 75454 74528 75486
rect 74208 75218 74250 75454
rect 74486 75218 74528 75454
rect 74208 75134 74528 75218
rect 74208 74898 74250 75134
rect 74486 74898 74528 75134
rect 74208 74866 74528 74898
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 66000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 66000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 66000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 66000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 86726 5133 86786 567291
rect 89568 561454 89888 561486
rect 89568 561218 89610 561454
rect 89846 561218 89888 561454
rect 89568 561134 89888 561218
rect 89568 560898 89610 561134
rect 89846 560898 89888 561134
rect 89568 560866 89888 560898
rect 89568 525454 89888 525486
rect 89568 525218 89610 525454
rect 89846 525218 89888 525454
rect 89568 525134 89888 525218
rect 89568 524898 89610 525134
rect 89846 524898 89888 525134
rect 89568 524866 89888 524898
rect 89568 489454 89888 489486
rect 89568 489218 89610 489454
rect 89846 489218 89888 489454
rect 89568 489134 89888 489218
rect 89568 488898 89610 489134
rect 89846 488898 89888 489134
rect 89568 488866 89888 488898
rect 89568 453454 89888 453486
rect 89568 453218 89610 453454
rect 89846 453218 89888 453454
rect 89568 453134 89888 453218
rect 89568 452898 89610 453134
rect 89846 452898 89888 453134
rect 89568 452866 89888 452898
rect 89568 417454 89888 417486
rect 89568 417218 89610 417454
rect 89846 417218 89888 417454
rect 89568 417134 89888 417218
rect 89568 416898 89610 417134
rect 89846 416898 89888 417134
rect 89568 416866 89888 416898
rect 89568 381454 89888 381486
rect 89568 381218 89610 381454
rect 89846 381218 89888 381454
rect 89568 381134 89888 381218
rect 89568 380898 89610 381134
rect 89846 380898 89888 381134
rect 89568 380866 89888 380898
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 89568 309454 89888 309486
rect 89568 309218 89610 309454
rect 89846 309218 89888 309454
rect 89568 309134 89888 309218
rect 89568 308898 89610 309134
rect 89846 308898 89888 309134
rect 89568 308866 89888 308898
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 89568 237454 89888 237486
rect 89568 237218 89610 237454
rect 89846 237218 89888 237454
rect 89568 237134 89888 237218
rect 89568 236898 89610 237134
rect 89846 236898 89888 237134
rect 89568 236866 89888 236898
rect 89568 201454 89888 201486
rect 89568 201218 89610 201454
rect 89846 201218 89888 201454
rect 89568 201134 89888 201218
rect 89568 200898 89610 201134
rect 89846 200898 89888 201134
rect 89568 200866 89888 200898
rect 89568 165454 89888 165486
rect 89568 165218 89610 165454
rect 89846 165218 89888 165454
rect 89568 165134 89888 165218
rect 89568 164898 89610 165134
rect 89846 164898 89888 165134
rect 89568 164866 89888 164898
rect 89568 129454 89888 129486
rect 89568 129218 89610 129454
rect 89846 129218 89888 129454
rect 89568 129134 89888 129218
rect 89568 128898 89610 129134
rect 89846 128898 89888 129134
rect 89568 128866 89888 128898
rect 89568 93454 89888 93486
rect 89568 93218 89610 93454
rect 89846 93218 89888 93454
rect 89568 93134 89888 93218
rect 89568 92898 89610 93134
rect 89846 92898 89888 93134
rect 89568 92866 89888 92898
rect 91794 57454 92414 66000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 86723 5132 86789 5133
rect 86723 5068 86724 5132
rect 86788 5068 86789 5132
rect 86723 5067 86789 5068
rect 91794 -1306 92414 20898
rect 93718 3501 93778 570691
rect 95514 570000 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 97763 570620 97829 570621
rect 97763 570556 97764 570620
rect 97828 570556 97829 570620
rect 97763 570555 97829 570556
rect 95514 61174 96134 66000
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 93715 3500 93781 3501
rect 93715 3436 93716 3500
rect 93780 3436 93781 3500
rect 93715 3435 93781 3436
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 -3226 96134 24618
rect 97766 3501 97826 570555
rect 99234 570000 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 106779 699820 106845 699821
rect 106779 699756 106780 699820
rect 106844 699756 106845 699820
rect 106779 699755 106845 699756
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 570000 103574 572058
rect 101995 567356 102061 567357
rect 101995 567292 101996 567356
rect 102060 567292 102061 567356
rect 101995 567291 102061 567292
rect 99234 64894 99854 66000
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 97763 3500 97829 3501
rect 97763 3436 97764 3500
rect 97828 3436 97829 3500
rect 97763 3435 97829 3436
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 28338
rect 101998 6493 102058 567291
rect 104928 543454 105248 543486
rect 104928 543218 104970 543454
rect 105206 543218 105248 543454
rect 104928 543134 105248 543218
rect 104928 542898 104970 543134
rect 105206 542898 105248 543134
rect 104928 542866 105248 542898
rect 104928 507454 105248 507486
rect 104928 507218 104970 507454
rect 105206 507218 105248 507454
rect 104928 507134 105248 507218
rect 104928 506898 104970 507134
rect 105206 506898 105248 507134
rect 104928 506866 105248 506898
rect 104928 471454 105248 471486
rect 104928 471218 104970 471454
rect 105206 471218 105248 471454
rect 104928 471134 105248 471218
rect 104928 470898 104970 471134
rect 105206 470898 105248 471134
rect 104928 470866 105248 470898
rect 104928 435454 105248 435486
rect 104928 435218 104970 435454
rect 105206 435218 105248 435454
rect 104928 435134 105248 435218
rect 104928 434898 104970 435134
rect 105206 434898 105248 435134
rect 104928 434866 105248 434898
rect 104928 399454 105248 399486
rect 104928 399218 104970 399454
rect 105206 399218 105248 399454
rect 104928 399134 105248 399218
rect 104928 398898 104970 399134
rect 105206 398898 105248 399134
rect 104928 398866 105248 398898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 104928 327454 105248 327486
rect 104928 327218 104970 327454
rect 105206 327218 105248 327454
rect 104928 327134 105248 327218
rect 104928 326898 104970 327134
rect 105206 326898 105248 327134
rect 104928 326866 105248 326898
rect 104928 291454 105248 291486
rect 104928 291218 104970 291454
rect 105206 291218 105248 291454
rect 104928 291134 105248 291218
rect 104928 290898 104970 291134
rect 105206 290898 105248 291134
rect 104928 290866 105248 290898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 104928 219454 105248 219486
rect 104928 219218 104970 219454
rect 105206 219218 105248 219454
rect 104928 219134 105248 219218
rect 104928 218898 104970 219134
rect 105206 218898 105248 219134
rect 104928 218866 105248 218898
rect 104928 183454 105248 183486
rect 104928 183218 104970 183454
rect 105206 183218 105248 183454
rect 104928 183134 105248 183218
rect 104928 182898 104970 183134
rect 105206 182898 105248 183134
rect 104928 182866 105248 182898
rect 104928 147454 105248 147486
rect 104928 147218 104970 147454
rect 105206 147218 105248 147454
rect 104928 147134 105248 147218
rect 104928 146898 104970 147134
rect 105206 146898 105248 147134
rect 104928 146866 105248 146898
rect 104928 111454 105248 111486
rect 104928 111218 104970 111454
rect 105206 111218 105248 111454
rect 104928 111134 105248 111218
rect 104928 110898 104970 111134
rect 105206 110898 105248 111134
rect 104928 110866 105248 110898
rect 104928 75454 105248 75486
rect 104928 75218 104970 75454
rect 105206 75218 105248 75454
rect 104928 75134 105248 75218
rect 104928 74898 104970 75134
rect 105206 74898 105248 75134
rect 104928 74866 105248 74898
rect 106782 67421 106842 699755
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 570000 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111563 570892 111629 570893
rect 111563 570828 111564 570892
rect 111628 570828 111629 570892
rect 111563 570827 111629 570828
rect 106779 67420 106845 67421
rect 106779 67356 106780 67420
rect 106844 67356 106845 67420
rect 106779 67355 106845 67356
rect 102954 32614 103574 66000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 101995 6492 102061 6493
rect 101995 6428 101996 6492
rect 102060 6428 102061 6492
rect 101995 6427 102061 6428
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 66000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 111566 3501 111626 570827
rect 113514 570000 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 570000 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 570000 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 570000 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 570000 132134 600618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 570000 135854 604338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 570000 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145603 570212 145669 570213
rect 145603 570148 145604 570212
rect 145668 570148 145669 570212
rect 145603 570147 145669 570148
rect 133643 567356 133709 567357
rect 133643 567292 133644 567356
rect 133708 567292 133709 567356
rect 133643 567291 133709 567292
rect 144683 567356 144749 567357
rect 144683 567292 144684 567356
rect 144748 567292 144749 567356
rect 144683 567291 144749 567292
rect 130883 566540 130949 566541
rect 130883 566476 130884 566540
rect 130948 566476 130949 566540
rect 130883 566475 130949 566476
rect 120288 561454 120608 561486
rect 120288 561218 120330 561454
rect 120566 561218 120608 561454
rect 120288 561134 120608 561218
rect 120288 560898 120330 561134
rect 120566 560898 120608 561134
rect 120288 560866 120608 560898
rect 120288 525454 120608 525486
rect 120288 525218 120330 525454
rect 120566 525218 120608 525454
rect 120288 525134 120608 525218
rect 120288 524898 120330 525134
rect 120566 524898 120608 525134
rect 120288 524866 120608 524898
rect 120288 489454 120608 489486
rect 120288 489218 120330 489454
rect 120566 489218 120608 489454
rect 120288 489134 120608 489218
rect 120288 488898 120330 489134
rect 120566 488898 120608 489134
rect 120288 488866 120608 488898
rect 120288 453454 120608 453486
rect 120288 453218 120330 453454
rect 120566 453218 120608 453454
rect 120288 453134 120608 453218
rect 120288 452898 120330 453134
rect 120566 452898 120608 453134
rect 120288 452866 120608 452898
rect 120288 417454 120608 417486
rect 120288 417218 120330 417454
rect 120566 417218 120608 417454
rect 120288 417134 120608 417218
rect 120288 416898 120330 417134
rect 120566 416898 120608 417134
rect 120288 416866 120608 416898
rect 120288 381454 120608 381486
rect 120288 381218 120330 381454
rect 120566 381218 120608 381454
rect 120288 381134 120608 381218
rect 120288 380898 120330 381134
rect 120566 380898 120608 381134
rect 120288 380866 120608 380898
rect 120288 345454 120608 345486
rect 120288 345218 120330 345454
rect 120566 345218 120608 345454
rect 120288 345134 120608 345218
rect 120288 344898 120330 345134
rect 120566 344898 120608 345134
rect 120288 344866 120608 344898
rect 120288 309454 120608 309486
rect 120288 309218 120330 309454
rect 120566 309218 120608 309454
rect 120288 309134 120608 309218
rect 120288 308898 120330 309134
rect 120566 308898 120608 309134
rect 120288 308866 120608 308898
rect 120288 273454 120608 273486
rect 120288 273218 120330 273454
rect 120566 273218 120608 273454
rect 120288 273134 120608 273218
rect 120288 272898 120330 273134
rect 120566 272898 120608 273134
rect 120288 272866 120608 272898
rect 120288 237454 120608 237486
rect 120288 237218 120330 237454
rect 120566 237218 120608 237454
rect 120288 237134 120608 237218
rect 120288 236898 120330 237134
rect 120566 236898 120608 237134
rect 120288 236866 120608 236898
rect 120288 201454 120608 201486
rect 120288 201218 120330 201454
rect 120566 201218 120608 201454
rect 120288 201134 120608 201218
rect 120288 200898 120330 201134
rect 120566 200898 120608 201134
rect 120288 200866 120608 200898
rect 120288 165454 120608 165486
rect 120288 165218 120330 165454
rect 120566 165218 120608 165454
rect 120288 165134 120608 165218
rect 120288 164898 120330 165134
rect 120566 164898 120608 165134
rect 120288 164866 120608 164898
rect 120288 129454 120608 129486
rect 120288 129218 120330 129454
rect 120566 129218 120608 129454
rect 120288 129134 120608 129218
rect 120288 128898 120330 129134
rect 120566 128898 120608 129134
rect 120288 128866 120608 128898
rect 120288 93454 120608 93486
rect 120288 93218 120330 93454
rect 120566 93218 120608 93454
rect 120288 93134 120608 93218
rect 120288 92898 120330 93134
rect 120566 92898 120608 93134
rect 120288 92866 120608 92898
rect 113514 43174 114134 66000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 111563 3500 111629 3501
rect 111563 3436 111564 3500
rect 111628 3436 111629 3500
rect 111563 3435 111629 3436
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 66000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 66000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 66000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 130886 3773 130946 566475
rect 131514 61174 132134 66000
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 130883 3772 130949 3773
rect 130883 3708 130884 3772
rect 130948 3708 130949 3772
rect 130883 3707 130949 3708
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 -3226 132134 24618
rect 133646 5541 133706 567291
rect 140635 566404 140701 566405
rect 140635 566340 140636 566404
rect 140700 566340 140701 566404
rect 140635 566339 140701 566340
rect 135648 543454 135968 543486
rect 135648 543218 135690 543454
rect 135926 543218 135968 543454
rect 135648 543134 135968 543218
rect 135648 542898 135690 543134
rect 135926 542898 135968 543134
rect 135648 542866 135968 542898
rect 135648 507454 135968 507486
rect 135648 507218 135690 507454
rect 135926 507218 135968 507454
rect 135648 507134 135968 507218
rect 135648 506898 135690 507134
rect 135926 506898 135968 507134
rect 135648 506866 135968 506898
rect 135648 471454 135968 471486
rect 135648 471218 135690 471454
rect 135926 471218 135968 471454
rect 135648 471134 135968 471218
rect 135648 470898 135690 471134
rect 135926 470898 135968 471134
rect 135648 470866 135968 470898
rect 135648 435454 135968 435486
rect 135648 435218 135690 435454
rect 135926 435218 135968 435454
rect 135648 435134 135968 435218
rect 135648 434898 135690 435134
rect 135926 434898 135968 435134
rect 135648 434866 135968 434898
rect 135648 399454 135968 399486
rect 135648 399218 135690 399454
rect 135926 399218 135968 399454
rect 135648 399134 135968 399218
rect 135648 398898 135690 399134
rect 135926 398898 135968 399134
rect 135648 398866 135968 398898
rect 135648 363454 135968 363486
rect 135648 363218 135690 363454
rect 135926 363218 135968 363454
rect 135648 363134 135968 363218
rect 135648 362898 135690 363134
rect 135926 362898 135968 363134
rect 135648 362866 135968 362898
rect 135648 327454 135968 327486
rect 135648 327218 135690 327454
rect 135926 327218 135968 327454
rect 135648 327134 135968 327218
rect 135648 326898 135690 327134
rect 135926 326898 135968 327134
rect 135648 326866 135968 326898
rect 135648 291454 135968 291486
rect 135648 291218 135690 291454
rect 135926 291218 135968 291454
rect 135648 291134 135968 291218
rect 135648 290898 135690 291134
rect 135926 290898 135968 291134
rect 135648 290866 135968 290898
rect 135648 255454 135968 255486
rect 135648 255218 135690 255454
rect 135926 255218 135968 255454
rect 135648 255134 135968 255218
rect 135648 254898 135690 255134
rect 135926 254898 135968 255134
rect 135648 254866 135968 254898
rect 135648 219454 135968 219486
rect 135648 219218 135690 219454
rect 135926 219218 135968 219454
rect 135648 219134 135968 219218
rect 135648 218898 135690 219134
rect 135926 218898 135968 219134
rect 135648 218866 135968 218898
rect 135648 183454 135968 183486
rect 135648 183218 135690 183454
rect 135926 183218 135968 183454
rect 135648 183134 135968 183218
rect 135648 182898 135690 183134
rect 135926 182898 135968 183134
rect 135648 182866 135968 182898
rect 135648 147454 135968 147486
rect 135648 147218 135690 147454
rect 135926 147218 135968 147454
rect 135648 147134 135968 147218
rect 135648 146898 135690 147134
rect 135926 146898 135968 147134
rect 135648 146866 135968 146898
rect 135648 111454 135968 111486
rect 135648 111218 135690 111454
rect 135926 111218 135968 111454
rect 135648 111134 135968 111218
rect 135648 110898 135690 111134
rect 135926 110898 135968 111134
rect 135648 110866 135968 110898
rect 135648 75454 135968 75486
rect 135648 75218 135690 75454
rect 135926 75218 135968 75454
rect 135648 75134 135968 75218
rect 135648 74898 135690 75134
rect 135926 74898 135968 75134
rect 135648 74866 135968 74898
rect 135234 64894 135854 66000
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 133643 5540 133709 5541
rect 133643 5476 133644 5540
rect 133708 5476 133709 5540
rect 133643 5475 133709 5476
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 66000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 140638 3773 140698 566339
rect 144686 5405 144746 567291
rect 144683 5404 144749 5405
rect 144683 5340 144684 5404
rect 144748 5340 144749 5404
rect 144683 5339 144749 5340
rect 145606 3773 145666 570147
rect 145794 570000 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 570000 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 152963 571300 153029 571301
rect 152963 571236 152964 571300
rect 153028 571236 153029 571300
rect 152963 571235 153029 571236
rect 151008 561454 151328 561486
rect 151008 561218 151050 561454
rect 151286 561218 151328 561454
rect 151008 561134 151328 561218
rect 151008 560898 151050 561134
rect 151286 560898 151328 561134
rect 151008 560866 151328 560898
rect 151008 525454 151328 525486
rect 151008 525218 151050 525454
rect 151286 525218 151328 525454
rect 151008 525134 151328 525218
rect 151008 524898 151050 525134
rect 151286 524898 151328 525134
rect 151008 524866 151328 524898
rect 151008 489454 151328 489486
rect 151008 489218 151050 489454
rect 151286 489218 151328 489454
rect 151008 489134 151328 489218
rect 151008 488898 151050 489134
rect 151286 488898 151328 489134
rect 151008 488866 151328 488898
rect 151008 453454 151328 453486
rect 151008 453218 151050 453454
rect 151286 453218 151328 453454
rect 151008 453134 151328 453218
rect 151008 452898 151050 453134
rect 151286 452898 151328 453134
rect 151008 452866 151328 452898
rect 151008 417454 151328 417486
rect 151008 417218 151050 417454
rect 151286 417218 151328 417454
rect 151008 417134 151328 417218
rect 151008 416898 151050 417134
rect 151286 416898 151328 417134
rect 151008 416866 151328 416898
rect 151008 381454 151328 381486
rect 151008 381218 151050 381454
rect 151286 381218 151328 381454
rect 151008 381134 151328 381218
rect 151008 380898 151050 381134
rect 151286 380898 151328 381134
rect 151008 380866 151328 380898
rect 151008 345454 151328 345486
rect 151008 345218 151050 345454
rect 151286 345218 151328 345454
rect 151008 345134 151328 345218
rect 151008 344898 151050 345134
rect 151286 344898 151328 345134
rect 151008 344866 151328 344898
rect 151008 309454 151328 309486
rect 151008 309218 151050 309454
rect 151286 309218 151328 309454
rect 151008 309134 151328 309218
rect 151008 308898 151050 309134
rect 151286 308898 151328 309134
rect 151008 308866 151328 308898
rect 151008 273454 151328 273486
rect 151008 273218 151050 273454
rect 151286 273218 151328 273454
rect 151008 273134 151328 273218
rect 151008 272898 151050 273134
rect 151286 272898 151328 273134
rect 151008 272866 151328 272898
rect 151008 237454 151328 237486
rect 151008 237218 151050 237454
rect 151286 237218 151328 237454
rect 151008 237134 151328 237218
rect 151008 236898 151050 237134
rect 151286 236898 151328 237134
rect 151008 236866 151328 236898
rect 151008 201454 151328 201486
rect 151008 201218 151050 201454
rect 151286 201218 151328 201454
rect 151008 201134 151328 201218
rect 151008 200898 151050 201134
rect 151286 200898 151328 201134
rect 151008 200866 151328 200898
rect 151008 165454 151328 165486
rect 151008 165218 151050 165454
rect 151286 165218 151328 165454
rect 151008 165134 151328 165218
rect 151008 164898 151050 165134
rect 151286 164898 151328 165134
rect 151008 164866 151328 164898
rect 151008 129454 151328 129486
rect 151008 129218 151050 129454
rect 151286 129218 151328 129454
rect 151008 129134 151328 129218
rect 151008 128898 151050 129134
rect 151286 128898 151328 129134
rect 151008 128866 151328 128898
rect 151008 93454 151328 93486
rect 151008 93218 151050 93454
rect 151286 93218 151328 93454
rect 151008 93134 151328 93218
rect 151008 92898 151050 93134
rect 151286 92898 151328 93134
rect 151008 92866 151328 92898
rect 145794 39454 146414 66000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 140635 3772 140701 3773
rect 140635 3708 140636 3772
rect 140700 3708 140701 3772
rect 140635 3707 140701 3708
rect 145603 3772 145669 3773
rect 145603 3708 145604 3772
rect 145668 3708 145669 3772
rect 145603 3707 145669 3708
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 66000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 152966 3773 153026 571235
rect 153234 570000 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156643 571028 156709 571029
rect 156643 570964 156644 571028
rect 156708 570964 156709 571028
rect 156643 570963 156709 570964
rect 155723 567356 155789 567357
rect 155723 567292 155724 567356
rect 155788 567292 155789 567356
rect 155723 567291 155789 567292
rect 153234 46894 153854 66000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 152963 3772 153029 3773
rect 152963 3708 152964 3772
rect 153028 3708 153029 3772
rect 152963 3707 153029 3708
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 10338
rect 155726 5133 155786 567291
rect 155723 5132 155789 5133
rect 155723 5068 155724 5132
rect 155788 5068 155789 5132
rect 155723 5067 155789 5068
rect 156646 3773 156706 570963
rect 156954 570000 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 161243 570348 161309 570349
rect 161243 570284 161244 570348
rect 161308 570284 161309 570348
rect 161243 570283 161309 570284
rect 156954 50614 157574 66000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156643 3772 156709 3773
rect 156643 3708 156644 3772
rect 156708 3708 156709 3772
rect 156643 3707 156709 3708
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 161246 3773 161306 570283
rect 163794 570000 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 570000 168134 600618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 168971 570484 169037 570485
rect 168971 570420 168972 570484
rect 169036 570420 169037 570484
rect 168971 570419 169037 570420
rect 164555 566676 164621 566677
rect 164555 566612 164556 566676
rect 164620 566612 164621 566676
rect 164555 566611 164621 566612
rect 163794 57454 164414 66000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 161243 3772 161309 3773
rect 161243 3708 161244 3772
rect 161308 3708 161309 3772
rect 161243 3707 161309 3708
rect 163794 -1306 164414 20898
rect 164558 3773 164618 566611
rect 166368 543454 166688 543486
rect 166368 543218 166410 543454
rect 166646 543218 166688 543454
rect 166368 543134 166688 543218
rect 166368 542898 166410 543134
rect 166646 542898 166688 543134
rect 166368 542866 166688 542898
rect 166368 507454 166688 507486
rect 166368 507218 166410 507454
rect 166646 507218 166688 507454
rect 166368 507134 166688 507218
rect 166368 506898 166410 507134
rect 166646 506898 166688 507134
rect 166368 506866 166688 506898
rect 166368 471454 166688 471486
rect 166368 471218 166410 471454
rect 166646 471218 166688 471454
rect 166368 471134 166688 471218
rect 166368 470898 166410 471134
rect 166646 470898 166688 471134
rect 166368 470866 166688 470898
rect 166368 435454 166688 435486
rect 166368 435218 166410 435454
rect 166646 435218 166688 435454
rect 166368 435134 166688 435218
rect 166368 434898 166410 435134
rect 166646 434898 166688 435134
rect 166368 434866 166688 434898
rect 166368 399454 166688 399486
rect 166368 399218 166410 399454
rect 166646 399218 166688 399454
rect 166368 399134 166688 399218
rect 166368 398898 166410 399134
rect 166646 398898 166688 399134
rect 166368 398866 166688 398898
rect 166368 363454 166688 363486
rect 166368 363218 166410 363454
rect 166646 363218 166688 363454
rect 166368 363134 166688 363218
rect 166368 362898 166410 363134
rect 166646 362898 166688 363134
rect 166368 362866 166688 362898
rect 166368 327454 166688 327486
rect 166368 327218 166410 327454
rect 166646 327218 166688 327454
rect 166368 327134 166688 327218
rect 166368 326898 166410 327134
rect 166646 326898 166688 327134
rect 166368 326866 166688 326898
rect 166368 291454 166688 291486
rect 166368 291218 166410 291454
rect 166646 291218 166688 291454
rect 166368 291134 166688 291218
rect 166368 290898 166410 291134
rect 166646 290898 166688 291134
rect 166368 290866 166688 290898
rect 166368 255454 166688 255486
rect 166368 255218 166410 255454
rect 166646 255218 166688 255454
rect 166368 255134 166688 255218
rect 166368 254898 166410 255134
rect 166646 254898 166688 255134
rect 166368 254866 166688 254898
rect 166368 219454 166688 219486
rect 166368 219218 166410 219454
rect 166646 219218 166688 219454
rect 166368 219134 166688 219218
rect 166368 218898 166410 219134
rect 166646 218898 166688 219134
rect 166368 218866 166688 218898
rect 166368 183454 166688 183486
rect 166368 183218 166410 183454
rect 166646 183218 166688 183454
rect 166368 183134 166688 183218
rect 166368 182898 166410 183134
rect 166646 182898 166688 183134
rect 166368 182866 166688 182898
rect 166368 147454 166688 147486
rect 166368 147218 166410 147454
rect 166646 147218 166688 147454
rect 166368 147134 166688 147218
rect 166368 146898 166410 147134
rect 166646 146898 166688 147134
rect 166368 146866 166688 146898
rect 166368 111454 166688 111486
rect 166368 111218 166410 111454
rect 166646 111218 166688 111454
rect 166368 111134 166688 111218
rect 166368 110898 166410 111134
rect 166646 110898 166688 111134
rect 166368 110866 166688 110898
rect 166368 75454 166688 75486
rect 166368 75218 166410 75454
rect 166646 75218 166688 75454
rect 166368 75134 166688 75218
rect 166368 74898 166410 75134
rect 166646 74898 166688 75134
rect 166368 74866 166688 74898
rect 167514 61174 168134 66000
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 164555 3772 164621 3773
rect 164555 3708 164556 3772
rect 164620 3708 164621 3772
rect 164555 3707 164621 3708
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 168974 4997 169034 570419
rect 171234 570000 171854 604338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 570000 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 175779 571164 175845 571165
rect 175779 571100 175780 571164
rect 175844 571100 175845 571164
rect 175779 571099 175845 571100
rect 170995 567356 171061 567357
rect 170995 567292 170996 567356
rect 171060 567292 171061 567356
rect 170995 567291 171061 567292
rect 170998 5133 171058 567291
rect 171234 64894 171854 66000
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 170995 5132 171061 5133
rect 170995 5068 170996 5132
rect 171060 5068 171061 5132
rect 170995 5067 171061 5068
rect 168971 4996 169037 4997
rect 168971 4932 168972 4996
rect 169036 4932 169037 4996
rect 168971 4931 169037 4932
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 66000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 175782 5269 175842 571099
rect 181794 570000 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 570000 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 570000 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 570000 193574 590058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 570000 200414 596898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 570000 204134 600618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 570000 207854 604338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 570000 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 570000 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 220675 570076 220741 570077
rect 220675 570012 220676 570076
rect 220740 570012 220741 570076
rect 220675 570011 220741 570012
rect 177987 568580 178053 568581
rect 177987 568516 177988 568580
rect 178052 568516 178053 568580
rect 177987 568515 178053 568516
rect 175779 5268 175845 5269
rect 175779 5204 175780 5268
rect 175844 5204 175845 5268
rect 175779 5203 175845 5204
rect 177990 3637 178050 568515
rect 210371 567356 210437 567357
rect 210371 567292 210372 567356
rect 210436 567292 210437 567356
rect 210371 567291 210437 567292
rect 210374 565997 210434 567291
rect 214419 567220 214485 567221
rect 214419 567156 214420 567220
rect 214484 567156 214485 567220
rect 214419 567155 214485 567156
rect 205403 565996 205469 565997
rect 205403 565932 205404 565996
rect 205468 565932 205469 565996
rect 205403 565931 205469 565932
rect 210371 565996 210437 565997
rect 210371 565932 210372 565996
rect 210436 565932 210437 565996
rect 210371 565931 210437 565932
rect 181728 561454 182048 561486
rect 181728 561218 181770 561454
rect 182006 561218 182048 561454
rect 181728 561134 182048 561218
rect 181728 560898 181770 561134
rect 182006 560898 182048 561134
rect 181728 560866 182048 560898
rect 197088 543454 197408 543486
rect 197088 543218 197130 543454
rect 197366 543218 197408 543454
rect 197088 543134 197408 543218
rect 197088 542898 197130 543134
rect 197366 542898 197408 543134
rect 197088 542866 197408 542898
rect 181728 525454 182048 525486
rect 181728 525218 181770 525454
rect 182006 525218 182048 525454
rect 181728 525134 182048 525218
rect 181728 524898 181770 525134
rect 182006 524898 182048 525134
rect 181728 524866 182048 524898
rect 197088 507454 197408 507486
rect 197088 507218 197130 507454
rect 197366 507218 197408 507454
rect 197088 507134 197408 507218
rect 197088 506898 197130 507134
rect 197366 506898 197408 507134
rect 197088 506866 197408 506898
rect 181728 489454 182048 489486
rect 181728 489218 181770 489454
rect 182006 489218 182048 489454
rect 181728 489134 182048 489218
rect 181728 488898 181770 489134
rect 182006 488898 182048 489134
rect 181728 488866 182048 488898
rect 197088 471454 197408 471486
rect 197088 471218 197130 471454
rect 197366 471218 197408 471454
rect 197088 471134 197408 471218
rect 197088 470898 197130 471134
rect 197366 470898 197408 471134
rect 197088 470866 197408 470898
rect 181728 453454 182048 453486
rect 181728 453218 181770 453454
rect 182006 453218 182048 453454
rect 181728 453134 182048 453218
rect 181728 452898 181770 453134
rect 182006 452898 182048 453134
rect 181728 452866 182048 452898
rect 197088 435454 197408 435486
rect 197088 435218 197130 435454
rect 197366 435218 197408 435454
rect 197088 435134 197408 435218
rect 197088 434898 197130 435134
rect 197366 434898 197408 435134
rect 197088 434866 197408 434898
rect 181728 417454 182048 417486
rect 181728 417218 181770 417454
rect 182006 417218 182048 417454
rect 181728 417134 182048 417218
rect 181728 416898 181770 417134
rect 182006 416898 182048 417134
rect 181728 416866 182048 416898
rect 197088 399454 197408 399486
rect 197088 399218 197130 399454
rect 197366 399218 197408 399454
rect 197088 399134 197408 399218
rect 197088 398898 197130 399134
rect 197366 398898 197408 399134
rect 197088 398866 197408 398898
rect 181728 381454 182048 381486
rect 181728 381218 181770 381454
rect 182006 381218 182048 381454
rect 181728 381134 182048 381218
rect 181728 380898 181770 381134
rect 182006 380898 182048 381134
rect 181728 380866 182048 380898
rect 197088 363454 197408 363486
rect 197088 363218 197130 363454
rect 197366 363218 197408 363454
rect 197088 363134 197408 363218
rect 197088 362898 197130 363134
rect 197366 362898 197408 363134
rect 197088 362866 197408 362898
rect 181728 345454 182048 345486
rect 181728 345218 181770 345454
rect 182006 345218 182048 345454
rect 181728 345134 182048 345218
rect 181728 344898 181770 345134
rect 182006 344898 182048 345134
rect 181728 344866 182048 344898
rect 197088 327454 197408 327486
rect 197088 327218 197130 327454
rect 197366 327218 197408 327454
rect 197088 327134 197408 327218
rect 197088 326898 197130 327134
rect 197366 326898 197408 327134
rect 197088 326866 197408 326898
rect 181728 309454 182048 309486
rect 181728 309218 181770 309454
rect 182006 309218 182048 309454
rect 181728 309134 182048 309218
rect 181728 308898 181770 309134
rect 182006 308898 182048 309134
rect 181728 308866 182048 308898
rect 197088 291454 197408 291486
rect 197088 291218 197130 291454
rect 197366 291218 197408 291454
rect 197088 291134 197408 291218
rect 197088 290898 197130 291134
rect 197366 290898 197408 291134
rect 197088 290866 197408 290898
rect 181728 273454 182048 273486
rect 181728 273218 181770 273454
rect 182006 273218 182048 273454
rect 181728 273134 182048 273218
rect 181728 272898 181770 273134
rect 182006 272898 182048 273134
rect 181728 272866 182048 272898
rect 197088 255454 197408 255486
rect 197088 255218 197130 255454
rect 197366 255218 197408 255454
rect 197088 255134 197408 255218
rect 197088 254898 197130 255134
rect 197366 254898 197408 255134
rect 197088 254866 197408 254898
rect 181728 237454 182048 237486
rect 181728 237218 181770 237454
rect 182006 237218 182048 237454
rect 181728 237134 182048 237218
rect 181728 236898 181770 237134
rect 182006 236898 182048 237134
rect 181728 236866 182048 236898
rect 197088 219454 197408 219486
rect 197088 219218 197130 219454
rect 197366 219218 197408 219454
rect 197088 219134 197408 219218
rect 197088 218898 197130 219134
rect 197366 218898 197408 219134
rect 197088 218866 197408 218898
rect 181728 201454 182048 201486
rect 181728 201218 181770 201454
rect 182006 201218 182048 201454
rect 181728 201134 182048 201218
rect 181728 200898 181770 201134
rect 182006 200898 182048 201134
rect 181728 200866 182048 200898
rect 197088 183454 197408 183486
rect 197088 183218 197130 183454
rect 197366 183218 197408 183454
rect 197088 183134 197408 183218
rect 197088 182898 197130 183134
rect 197366 182898 197408 183134
rect 197088 182866 197408 182898
rect 181728 165454 182048 165486
rect 181728 165218 181770 165454
rect 182006 165218 182048 165454
rect 181728 165134 182048 165218
rect 181728 164898 181770 165134
rect 182006 164898 182048 165134
rect 181728 164866 182048 164898
rect 197088 147454 197408 147486
rect 197088 147218 197130 147454
rect 197366 147218 197408 147454
rect 197088 147134 197408 147218
rect 197088 146898 197130 147134
rect 197366 146898 197408 147134
rect 197088 146866 197408 146898
rect 181728 129454 182048 129486
rect 181728 129218 181770 129454
rect 182006 129218 182048 129454
rect 181728 129134 182048 129218
rect 181728 128898 181770 129134
rect 182006 128898 182048 129134
rect 181728 128866 182048 128898
rect 197088 111454 197408 111486
rect 197088 111218 197130 111454
rect 197366 111218 197408 111454
rect 197088 111134 197408 111218
rect 197088 110898 197130 111134
rect 197366 110898 197408 111134
rect 197088 110866 197408 110898
rect 181728 93454 182048 93486
rect 181728 93218 181770 93454
rect 182006 93218 182048 93454
rect 181728 93134 182048 93218
rect 181728 92898 181770 93134
rect 182006 92898 182048 93134
rect 181728 92866 182048 92898
rect 197088 75454 197408 75486
rect 197088 75218 197130 75454
rect 197366 75218 197408 75454
rect 197088 75134 197408 75218
rect 197088 74898 197130 75134
rect 197366 74898 197408 75134
rect 197088 74866 197408 74898
rect 181794 39454 182414 66000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 177987 3636 178053 3637
rect 177987 3572 177988 3636
rect 178052 3572 178053 3636
rect 177987 3571 178053 3572
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 66000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 66000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 66000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 66000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 66000
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 205406 3637 205466 565931
rect 212448 561454 212768 561486
rect 212448 561218 212490 561454
rect 212726 561218 212768 561454
rect 212448 561134 212768 561218
rect 212448 560898 212490 561134
rect 212726 560898 212768 561134
rect 212448 560866 212768 560898
rect 212448 525454 212768 525486
rect 212448 525218 212490 525454
rect 212726 525218 212768 525454
rect 212448 525134 212768 525218
rect 212448 524898 212490 525134
rect 212726 524898 212768 525134
rect 212448 524866 212768 524898
rect 212448 489454 212768 489486
rect 212448 489218 212490 489454
rect 212726 489218 212768 489454
rect 212448 489134 212768 489218
rect 212448 488898 212490 489134
rect 212726 488898 212768 489134
rect 212448 488866 212768 488898
rect 212448 453454 212768 453486
rect 212448 453218 212490 453454
rect 212726 453218 212768 453454
rect 212448 453134 212768 453218
rect 212448 452898 212490 453134
rect 212726 452898 212768 453134
rect 212448 452866 212768 452898
rect 212448 417454 212768 417486
rect 212448 417218 212490 417454
rect 212726 417218 212768 417454
rect 212448 417134 212768 417218
rect 212448 416898 212490 417134
rect 212726 416898 212768 417134
rect 212448 416866 212768 416898
rect 212448 381454 212768 381486
rect 212448 381218 212490 381454
rect 212726 381218 212768 381454
rect 212448 381134 212768 381218
rect 212448 380898 212490 381134
rect 212726 380898 212768 381134
rect 212448 380866 212768 380898
rect 212448 345454 212768 345486
rect 212448 345218 212490 345454
rect 212726 345218 212768 345454
rect 212448 345134 212768 345218
rect 212448 344898 212490 345134
rect 212726 344898 212768 345134
rect 212448 344866 212768 344898
rect 212448 309454 212768 309486
rect 212448 309218 212490 309454
rect 212726 309218 212768 309454
rect 212448 309134 212768 309218
rect 212448 308898 212490 309134
rect 212726 308898 212768 309134
rect 212448 308866 212768 308898
rect 212448 273454 212768 273486
rect 212448 273218 212490 273454
rect 212726 273218 212768 273454
rect 212448 273134 212768 273218
rect 212448 272898 212490 273134
rect 212726 272898 212768 273134
rect 212448 272866 212768 272898
rect 212448 237454 212768 237486
rect 212448 237218 212490 237454
rect 212726 237218 212768 237454
rect 212448 237134 212768 237218
rect 212448 236898 212490 237134
rect 212726 236898 212768 237134
rect 212448 236866 212768 236898
rect 212448 201454 212768 201486
rect 212448 201218 212490 201454
rect 212726 201218 212768 201454
rect 212448 201134 212768 201218
rect 212448 200898 212490 201134
rect 212726 200898 212768 201134
rect 212448 200866 212768 200898
rect 212448 165454 212768 165486
rect 212448 165218 212490 165454
rect 212726 165218 212768 165454
rect 212448 165134 212768 165218
rect 212448 164898 212490 165134
rect 212726 164898 212768 165134
rect 212448 164866 212768 164898
rect 212448 129454 212768 129486
rect 212448 129218 212490 129454
rect 212726 129218 212768 129454
rect 212448 129134 212768 129218
rect 212448 128898 212490 129134
rect 212726 128898 212768 129134
rect 212448 128866 212768 128898
rect 212448 93454 212768 93486
rect 212448 93218 212490 93454
rect 212726 93218 212768 93454
rect 212448 93134 212768 93218
rect 212448 92898 212490 93134
rect 212726 92898 212768 93134
rect 212448 92866 212768 92898
rect 207234 64894 207854 66000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 205403 3636 205469 3637
rect 205403 3572 205404 3636
rect 205468 3572 205469 3636
rect 205403 3571 205469 3572
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 66000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 214422 3637 214482 567155
rect 217794 39454 218414 66000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 214419 3636 214485 3637
rect 214419 3572 214420 3636
rect 214484 3572 214485 3636
rect 214419 3571 214485 3572
rect 217794 3454 218414 38898
rect 220678 3637 220738 570011
rect 221514 570000 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 570000 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 234659 699820 234725 699821
rect 234659 699756 234660 699820
rect 234724 699756 234725 699820
rect 234659 699755 234725 699756
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 227483 571028 227549 571029
rect 227483 570964 227484 571028
rect 227548 570964 227549 571028
rect 227483 570963 227549 570964
rect 221514 43174 222134 66000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 220675 3636 220741 3637
rect 220675 3572 220676 3636
rect 220740 3572 220741 3636
rect 220675 3571 220741 3572
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 66000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 227486 3637 227546 570963
rect 228954 570000 229574 590058
rect 227808 543454 228128 543486
rect 227808 543218 227850 543454
rect 228086 543218 228128 543454
rect 227808 543134 228128 543218
rect 227808 542898 227850 543134
rect 228086 542898 228128 543134
rect 227808 542866 228128 542898
rect 227808 507454 228128 507486
rect 227808 507218 227850 507454
rect 228086 507218 228128 507454
rect 227808 507134 228128 507218
rect 227808 506898 227850 507134
rect 228086 506898 228128 507134
rect 227808 506866 228128 506898
rect 227808 471454 228128 471486
rect 227808 471218 227850 471454
rect 228086 471218 228128 471454
rect 227808 471134 228128 471218
rect 227808 470898 227850 471134
rect 228086 470898 228128 471134
rect 227808 470866 228128 470898
rect 227808 435454 228128 435486
rect 227808 435218 227850 435454
rect 228086 435218 228128 435454
rect 227808 435134 228128 435218
rect 227808 434898 227850 435134
rect 228086 434898 228128 435134
rect 227808 434866 228128 434898
rect 227808 399454 228128 399486
rect 227808 399218 227850 399454
rect 228086 399218 228128 399454
rect 227808 399134 228128 399218
rect 227808 398898 227850 399134
rect 228086 398898 228128 399134
rect 227808 398866 228128 398898
rect 227808 363454 228128 363486
rect 227808 363218 227850 363454
rect 228086 363218 228128 363454
rect 227808 363134 228128 363218
rect 227808 362898 227850 363134
rect 228086 362898 228128 363134
rect 227808 362866 228128 362898
rect 227808 327454 228128 327486
rect 227808 327218 227850 327454
rect 228086 327218 228128 327454
rect 227808 327134 228128 327218
rect 227808 326898 227850 327134
rect 228086 326898 228128 327134
rect 227808 326866 228128 326898
rect 227808 291454 228128 291486
rect 227808 291218 227850 291454
rect 228086 291218 228128 291454
rect 227808 291134 228128 291218
rect 227808 290898 227850 291134
rect 228086 290898 228128 291134
rect 227808 290866 228128 290898
rect 227808 255454 228128 255486
rect 227808 255218 227850 255454
rect 228086 255218 228128 255454
rect 227808 255134 228128 255218
rect 227808 254898 227850 255134
rect 228086 254898 228128 255134
rect 227808 254866 228128 254898
rect 227808 219454 228128 219486
rect 227808 219218 227850 219454
rect 228086 219218 228128 219454
rect 227808 219134 228128 219218
rect 227808 218898 227850 219134
rect 228086 218898 228128 219134
rect 227808 218866 228128 218898
rect 227808 183454 228128 183486
rect 227808 183218 227850 183454
rect 228086 183218 228128 183454
rect 227808 183134 228128 183218
rect 227808 182898 227850 183134
rect 228086 182898 228128 183134
rect 227808 182866 228128 182898
rect 227808 147454 228128 147486
rect 227808 147218 227850 147454
rect 228086 147218 228128 147454
rect 227808 147134 228128 147218
rect 227808 146898 227850 147134
rect 228086 146898 228128 147134
rect 227808 146866 228128 146898
rect 227808 111454 228128 111486
rect 227808 111218 227850 111454
rect 228086 111218 228128 111454
rect 227808 111134 228128 111218
rect 227808 110898 227850 111134
rect 228086 110898 228128 111134
rect 227808 110866 228128 110898
rect 227808 75454 228128 75486
rect 227808 75218 227850 75454
rect 228086 75218 228128 75454
rect 227808 75134 228128 75218
rect 227808 74898 227850 75134
rect 228086 74898 228128 75134
rect 227808 74866 228128 74898
rect 234662 67285 234722 699755
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 570000 236414 596898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 570000 240134 600618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 570000 243854 604338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 570000 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 570000 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 570000 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 570000 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 570000 265574 590058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 570000 272414 596898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 570000 276134 600618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 570000 279854 604338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 570000 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 570000 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 570000 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 570000 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 570000 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 570000 308414 596898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 570000 312134 600618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 570000 315854 604338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 570000 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 570000 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 570000 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 570000 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 570000 337574 590058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 570000 344414 596898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 346899 570892 346965 570893
rect 346899 570828 346900 570892
rect 346964 570828 346965 570892
rect 346899 570827 346965 570828
rect 244227 567356 244293 567357
rect 244227 567292 244228 567356
rect 244292 567292 244293 567356
rect 244227 567291 244293 567292
rect 270539 567356 270605 567357
rect 270539 567292 270540 567356
rect 270604 567292 270605 567356
rect 270539 567291 270605 567292
rect 281579 567356 281645 567357
rect 281579 567292 281580 567356
rect 281644 567292 281645 567356
rect 281579 567291 281645 567292
rect 328499 567356 328565 567357
rect 328499 567292 328500 567356
rect 328564 567292 328565 567356
rect 328499 567291 328565 567292
rect 345059 567356 345125 567357
rect 345059 567292 345060 567356
rect 345124 567292 345125 567356
rect 345059 567291 345125 567292
rect 243168 561454 243488 561486
rect 243168 561218 243210 561454
rect 243446 561218 243488 561454
rect 243168 561134 243488 561218
rect 243168 560898 243210 561134
rect 243446 560898 243488 561134
rect 243168 560866 243488 560898
rect 243168 525454 243488 525486
rect 243168 525218 243210 525454
rect 243446 525218 243488 525454
rect 243168 525134 243488 525218
rect 243168 524898 243210 525134
rect 243446 524898 243488 525134
rect 243168 524866 243488 524898
rect 243168 489454 243488 489486
rect 243168 489218 243210 489454
rect 243446 489218 243488 489454
rect 243168 489134 243488 489218
rect 243168 488898 243210 489134
rect 243446 488898 243488 489134
rect 243168 488866 243488 488898
rect 243168 453454 243488 453486
rect 243168 453218 243210 453454
rect 243446 453218 243488 453454
rect 243168 453134 243488 453218
rect 243168 452898 243210 453134
rect 243446 452898 243488 453134
rect 243168 452866 243488 452898
rect 243168 417454 243488 417486
rect 243168 417218 243210 417454
rect 243446 417218 243488 417454
rect 243168 417134 243488 417218
rect 243168 416898 243210 417134
rect 243446 416898 243488 417134
rect 243168 416866 243488 416898
rect 243168 381454 243488 381486
rect 243168 381218 243210 381454
rect 243446 381218 243488 381454
rect 243168 381134 243488 381218
rect 243168 380898 243210 381134
rect 243446 380898 243488 381134
rect 243168 380866 243488 380898
rect 243168 345454 243488 345486
rect 243168 345218 243210 345454
rect 243446 345218 243488 345454
rect 243168 345134 243488 345218
rect 243168 344898 243210 345134
rect 243446 344898 243488 345134
rect 243168 344866 243488 344898
rect 243168 309454 243488 309486
rect 243168 309218 243210 309454
rect 243446 309218 243488 309454
rect 243168 309134 243488 309218
rect 243168 308898 243210 309134
rect 243446 308898 243488 309134
rect 243168 308866 243488 308898
rect 243168 273454 243488 273486
rect 243168 273218 243210 273454
rect 243446 273218 243488 273454
rect 243168 273134 243488 273218
rect 243168 272898 243210 273134
rect 243446 272898 243488 273134
rect 243168 272866 243488 272898
rect 243168 237454 243488 237486
rect 243168 237218 243210 237454
rect 243446 237218 243488 237454
rect 243168 237134 243488 237218
rect 243168 236898 243210 237134
rect 243446 236898 243488 237134
rect 243168 236866 243488 236898
rect 243168 201454 243488 201486
rect 243168 201218 243210 201454
rect 243446 201218 243488 201454
rect 243168 201134 243488 201218
rect 243168 200898 243210 201134
rect 243446 200898 243488 201134
rect 243168 200866 243488 200898
rect 243168 165454 243488 165486
rect 243168 165218 243210 165454
rect 243446 165218 243488 165454
rect 243168 165134 243488 165218
rect 243168 164898 243210 165134
rect 243446 164898 243488 165134
rect 243168 164866 243488 164898
rect 243168 129454 243488 129486
rect 243168 129218 243210 129454
rect 243446 129218 243488 129454
rect 243168 129134 243488 129218
rect 243168 128898 243210 129134
rect 243446 128898 243488 129134
rect 243168 128866 243488 128898
rect 243168 93454 243488 93486
rect 243168 93218 243210 93454
rect 243446 93218 243488 93454
rect 243168 93134 243488 93218
rect 243168 92898 243210 93134
rect 243446 92898 243488 93134
rect 243168 92866 243488 92898
rect 234659 67284 234725 67285
rect 234659 67220 234660 67284
rect 234724 67220 234725 67284
rect 234659 67219 234725 67220
rect 228954 50614 229574 66000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 227483 3636 227549 3637
rect 227483 3572 227484 3636
rect 227548 3572 227549 3636
rect 227483 3571 227549 3572
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 66000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 66000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 66000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 244230 5949 244290 567291
rect 258528 543454 258848 543486
rect 258528 543218 258570 543454
rect 258806 543218 258848 543454
rect 258528 543134 258848 543218
rect 258528 542898 258570 543134
rect 258806 542898 258848 543134
rect 258528 542866 258848 542898
rect 258528 507454 258848 507486
rect 258528 507218 258570 507454
rect 258806 507218 258848 507454
rect 258528 507134 258848 507218
rect 258528 506898 258570 507134
rect 258806 506898 258848 507134
rect 258528 506866 258848 506898
rect 258528 471454 258848 471486
rect 258528 471218 258570 471454
rect 258806 471218 258848 471454
rect 258528 471134 258848 471218
rect 258528 470898 258570 471134
rect 258806 470898 258848 471134
rect 258528 470866 258848 470898
rect 258528 435454 258848 435486
rect 258528 435218 258570 435454
rect 258806 435218 258848 435454
rect 258528 435134 258848 435218
rect 258528 434898 258570 435134
rect 258806 434898 258848 435134
rect 258528 434866 258848 434898
rect 258528 399454 258848 399486
rect 258528 399218 258570 399454
rect 258806 399218 258848 399454
rect 258528 399134 258848 399218
rect 258528 398898 258570 399134
rect 258806 398898 258848 399134
rect 258528 398866 258848 398898
rect 258528 363454 258848 363486
rect 258528 363218 258570 363454
rect 258806 363218 258848 363454
rect 258528 363134 258848 363218
rect 258528 362898 258570 363134
rect 258806 362898 258848 363134
rect 258528 362866 258848 362898
rect 258528 327454 258848 327486
rect 258528 327218 258570 327454
rect 258806 327218 258848 327454
rect 258528 327134 258848 327218
rect 258528 326898 258570 327134
rect 258806 326898 258848 327134
rect 258528 326866 258848 326898
rect 258528 291454 258848 291486
rect 258528 291218 258570 291454
rect 258806 291218 258848 291454
rect 258528 291134 258848 291218
rect 258528 290898 258570 291134
rect 258806 290898 258848 291134
rect 258528 290866 258848 290898
rect 258528 255454 258848 255486
rect 258528 255218 258570 255454
rect 258806 255218 258848 255454
rect 258528 255134 258848 255218
rect 258528 254898 258570 255134
rect 258806 254898 258848 255134
rect 258528 254866 258848 254898
rect 258528 219454 258848 219486
rect 258528 219218 258570 219454
rect 258806 219218 258848 219454
rect 258528 219134 258848 219218
rect 258528 218898 258570 219134
rect 258806 218898 258848 219134
rect 258528 218866 258848 218898
rect 258528 183454 258848 183486
rect 258528 183218 258570 183454
rect 258806 183218 258848 183454
rect 258528 183134 258848 183218
rect 258528 182898 258570 183134
rect 258806 182898 258848 183134
rect 258528 182866 258848 182898
rect 258528 147454 258848 147486
rect 258528 147218 258570 147454
rect 258806 147218 258848 147454
rect 258528 147134 258848 147218
rect 258528 146898 258570 147134
rect 258806 146898 258848 147134
rect 258528 146866 258848 146898
rect 258528 111454 258848 111486
rect 258528 111218 258570 111454
rect 258806 111218 258848 111454
rect 258528 111134 258848 111218
rect 258528 110898 258570 111134
rect 258806 110898 258848 111134
rect 258528 110866 258848 110898
rect 258528 75454 258848 75486
rect 258528 75218 258570 75454
rect 258806 75218 258848 75454
rect 258528 75134 258848 75218
rect 258528 74898 258570 75134
rect 258806 74898 258848 75134
rect 258528 74866 258848 74898
rect 246954 32614 247574 66000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 244227 5948 244293 5949
rect 244227 5884 244228 5948
rect 244292 5884 244293 5948
rect 244227 5883 244293 5884
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 66000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 66000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 66000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 66000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 270542 5269 270602 567291
rect 273888 561454 274208 561486
rect 273888 561218 273930 561454
rect 274166 561218 274208 561454
rect 273888 561134 274208 561218
rect 273888 560898 273930 561134
rect 274166 560898 274208 561134
rect 273888 560866 274208 560898
rect 273888 525454 274208 525486
rect 273888 525218 273930 525454
rect 274166 525218 274208 525454
rect 273888 525134 274208 525218
rect 273888 524898 273930 525134
rect 274166 524898 274208 525134
rect 273888 524866 274208 524898
rect 273888 489454 274208 489486
rect 273888 489218 273930 489454
rect 274166 489218 274208 489454
rect 273888 489134 274208 489218
rect 273888 488898 273930 489134
rect 274166 488898 274208 489134
rect 273888 488866 274208 488898
rect 273888 453454 274208 453486
rect 273888 453218 273930 453454
rect 274166 453218 274208 453454
rect 273888 453134 274208 453218
rect 273888 452898 273930 453134
rect 274166 452898 274208 453134
rect 273888 452866 274208 452898
rect 273888 417454 274208 417486
rect 273888 417218 273930 417454
rect 274166 417218 274208 417454
rect 273888 417134 274208 417218
rect 273888 416898 273930 417134
rect 274166 416898 274208 417134
rect 273888 416866 274208 416898
rect 273888 381454 274208 381486
rect 273888 381218 273930 381454
rect 274166 381218 274208 381454
rect 273888 381134 274208 381218
rect 273888 380898 273930 381134
rect 274166 380898 274208 381134
rect 273888 380866 274208 380898
rect 273888 345454 274208 345486
rect 273888 345218 273930 345454
rect 274166 345218 274208 345454
rect 273888 345134 274208 345218
rect 273888 344898 273930 345134
rect 274166 344898 274208 345134
rect 273888 344866 274208 344898
rect 273888 309454 274208 309486
rect 273888 309218 273930 309454
rect 274166 309218 274208 309454
rect 273888 309134 274208 309218
rect 273888 308898 273930 309134
rect 274166 308898 274208 309134
rect 273888 308866 274208 308898
rect 273888 273454 274208 273486
rect 273888 273218 273930 273454
rect 274166 273218 274208 273454
rect 273888 273134 274208 273218
rect 273888 272898 273930 273134
rect 274166 272898 274208 273134
rect 273888 272866 274208 272898
rect 273888 237454 274208 237486
rect 273888 237218 273930 237454
rect 274166 237218 274208 237454
rect 273888 237134 274208 237218
rect 273888 236898 273930 237134
rect 274166 236898 274208 237134
rect 273888 236866 274208 236898
rect 273888 201454 274208 201486
rect 273888 201218 273930 201454
rect 274166 201218 274208 201454
rect 273888 201134 274208 201218
rect 273888 200898 273930 201134
rect 274166 200898 274208 201134
rect 273888 200866 274208 200898
rect 273888 165454 274208 165486
rect 273888 165218 273930 165454
rect 274166 165218 274208 165454
rect 273888 165134 274208 165218
rect 273888 164898 273930 165134
rect 274166 164898 274208 165134
rect 273888 164866 274208 164898
rect 273888 129454 274208 129486
rect 273888 129218 273930 129454
rect 274166 129218 274208 129454
rect 273888 129134 274208 129218
rect 273888 128898 273930 129134
rect 274166 128898 274208 129134
rect 273888 128866 274208 128898
rect 273888 93454 274208 93486
rect 273888 93218 273930 93454
rect 274166 93218 274208 93454
rect 273888 93134 274208 93218
rect 273888 92898 273930 93134
rect 274166 92898 274208 93134
rect 273888 92866 274208 92898
rect 271794 57454 272414 66000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 270539 5268 270605 5269
rect 270539 5204 270540 5268
rect 270604 5204 270605 5268
rect 270539 5203 270605 5204
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 66000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 66000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 281582 6085 281642 567291
rect 328502 566541 328562 567291
rect 328499 566540 328565 566541
rect 328499 566476 328500 566540
rect 328564 566476 328565 566540
rect 328499 566475 328565 566476
rect 304608 561454 304928 561486
rect 304608 561218 304650 561454
rect 304886 561218 304928 561454
rect 304608 561134 304928 561218
rect 304608 560898 304650 561134
rect 304886 560898 304928 561134
rect 304608 560866 304928 560898
rect 335328 561454 335648 561486
rect 335328 561218 335370 561454
rect 335606 561218 335648 561454
rect 335328 561134 335648 561218
rect 335328 560898 335370 561134
rect 335606 560898 335648 561134
rect 335328 560866 335648 560898
rect 289248 543454 289568 543486
rect 289248 543218 289290 543454
rect 289526 543218 289568 543454
rect 289248 543134 289568 543218
rect 289248 542898 289290 543134
rect 289526 542898 289568 543134
rect 289248 542866 289568 542898
rect 319968 543454 320288 543486
rect 319968 543218 320010 543454
rect 320246 543218 320288 543454
rect 319968 543134 320288 543218
rect 319968 542898 320010 543134
rect 320246 542898 320288 543134
rect 319968 542866 320288 542898
rect 304608 525454 304928 525486
rect 304608 525218 304650 525454
rect 304886 525218 304928 525454
rect 304608 525134 304928 525218
rect 304608 524898 304650 525134
rect 304886 524898 304928 525134
rect 304608 524866 304928 524898
rect 335328 525454 335648 525486
rect 335328 525218 335370 525454
rect 335606 525218 335648 525454
rect 335328 525134 335648 525218
rect 335328 524898 335370 525134
rect 335606 524898 335648 525134
rect 335328 524866 335648 524898
rect 289248 507454 289568 507486
rect 289248 507218 289290 507454
rect 289526 507218 289568 507454
rect 289248 507134 289568 507218
rect 289248 506898 289290 507134
rect 289526 506898 289568 507134
rect 289248 506866 289568 506898
rect 319968 507454 320288 507486
rect 319968 507218 320010 507454
rect 320246 507218 320288 507454
rect 319968 507134 320288 507218
rect 319968 506898 320010 507134
rect 320246 506898 320288 507134
rect 319968 506866 320288 506898
rect 304608 489454 304928 489486
rect 304608 489218 304650 489454
rect 304886 489218 304928 489454
rect 304608 489134 304928 489218
rect 304608 488898 304650 489134
rect 304886 488898 304928 489134
rect 304608 488866 304928 488898
rect 335328 489454 335648 489486
rect 335328 489218 335370 489454
rect 335606 489218 335648 489454
rect 335328 489134 335648 489218
rect 335328 488898 335370 489134
rect 335606 488898 335648 489134
rect 335328 488866 335648 488898
rect 289248 471454 289568 471486
rect 289248 471218 289290 471454
rect 289526 471218 289568 471454
rect 289248 471134 289568 471218
rect 289248 470898 289290 471134
rect 289526 470898 289568 471134
rect 289248 470866 289568 470898
rect 319968 471454 320288 471486
rect 319968 471218 320010 471454
rect 320246 471218 320288 471454
rect 319968 471134 320288 471218
rect 319968 470898 320010 471134
rect 320246 470898 320288 471134
rect 319968 470866 320288 470898
rect 304608 453454 304928 453486
rect 304608 453218 304650 453454
rect 304886 453218 304928 453454
rect 304608 453134 304928 453218
rect 304608 452898 304650 453134
rect 304886 452898 304928 453134
rect 304608 452866 304928 452898
rect 335328 453454 335648 453486
rect 335328 453218 335370 453454
rect 335606 453218 335648 453454
rect 335328 453134 335648 453218
rect 335328 452898 335370 453134
rect 335606 452898 335648 453134
rect 335328 452866 335648 452898
rect 289248 435454 289568 435486
rect 289248 435218 289290 435454
rect 289526 435218 289568 435454
rect 289248 435134 289568 435218
rect 289248 434898 289290 435134
rect 289526 434898 289568 435134
rect 289248 434866 289568 434898
rect 319968 435454 320288 435486
rect 319968 435218 320010 435454
rect 320246 435218 320288 435454
rect 319968 435134 320288 435218
rect 319968 434898 320010 435134
rect 320246 434898 320288 435134
rect 319968 434866 320288 434898
rect 304608 417454 304928 417486
rect 304608 417218 304650 417454
rect 304886 417218 304928 417454
rect 304608 417134 304928 417218
rect 304608 416898 304650 417134
rect 304886 416898 304928 417134
rect 304608 416866 304928 416898
rect 335328 417454 335648 417486
rect 335328 417218 335370 417454
rect 335606 417218 335648 417454
rect 335328 417134 335648 417218
rect 335328 416898 335370 417134
rect 335606 416898 335648 417134
rect 335328 416866 335648 416898
rect 289248 399454 289568 399486
rect 289248 399218 289290 399454
rect 289526 399218 289568 399454
rect 289248 399134 289568 399218
rect 289248 398898 289290 399134
rect 289526 398898 289568 399134
rect 289248 398866 289568 398898
rect 319968 399454 320288 399486
rect 319968 399218 320010 399454
rect 320246 399218 320288 399454
rect 319968 399134 320288 399218
rect 319968 398898 320010 399134
rect 320246 398898 320288 399134
rect 319968 398866 320288 398898
rect 304608 381454 304928 381486
rect 304608 381218 304650 381454
rect 304886 381218 304928 381454
rect 304608 381134 304928 381218
rect 304608 380898 304650 381134
rect 304886 380898 304928 381134
rect 304608 380866 304928 380898
rect 335328 381454 335648 381486
rect 335328 381218 335370 381454
rect 335606 381218 335648 381454
rect 335328 381134 335648 381218
rect 335328 380898 335370 381134
rect 335606 380898 335648 381134
rect 335328 380866 335648 380898
rect 289248 363454 289568 363486
rect 289248 363218 289290 363454
rect 289526 363218 289568 363454
rect 289248 363134 289568 363218
rect 289248 362898 289290 363134
rect 289526 362898 289568 363134
rect 289248 362866 289568 362898
rect 319968 363454 320288 363486
rect 319968 363218 320010 363454
rect 320246 363218 320288 363454
rect 319968 363134 320288 363218
rect 319968 362898 320010 363134
rect 320246 362898 320288 363134
rect 319968 362866 320288 362898
rect 304608 345454 304928 345486
rect 304608 345218 304650 345454
rect 304886 345218 304928 345454
rect 304608 345134 304928 345218
rect 304608 344898 304650 345134
rect 304886 344898 304928 345134
rect 304608 344866 304928 344898
rect 335328 345454 335648 345486
rect 335328 345218 335370 345454
rect 335606 345218 335648 345454
rect 335328 345134 335648 345218
rect 335328 344898 335370 345134
rect 335606 344898 335648 345134
rect 335328 344866 335648 344898
rect 289248 327454 289568 327486
rect 289248 327218 289290 327454
rect 289526 327218 289568 327454
rect 289248 327134 289568 327218
rect 289248 326898 289290 327134
rect 289526 326898 289568 327134
rect 289248 326866 289568 326898
rect 319968 327454 320288 327486
rect 319968 327218 320010 327454
rect 320246 327218 320288 327454
rect 319968 327134 320288 327218
rect 319968 326898 320010 327134
rect 320246 326898 320288 327134
rect 319968 326866 320288 326898
rect 304608 309454 304928 309486
rect 304608 309218 304650 309454
rect 304886 309218 304928 309454
rect 304608 309134 304928 309218
rect 304608 308898 304650 309134
rect 304886 308898 304928 309134
rect 304608 308866 304928 308898
rect 335328 309454 335648 309486
rect 335328 309218 335370 309454
rect 335606 309218 335648 309454
rect 335328 309134 335648 309218
rect 335328 308898 335370 309134
rect 335606 308898 335648 309134
rect 335328 308866 335648 308898
rect 289248 291454 289568 291486
rect 289248 291218 289290 291454
rect 289526 291218 289568 291454
rect 289248 291134 289568 291218
rect 289248 290898 289290 291134
rect 289526 290898 289568 291134
rect 289248 290866 289568 290898
rect 319968 291454 320288 291486
rect 319968 291218 320010 291454
rect 320246 291218 320288 291454
rect 319968 291134 320288 291218
rect 319968 290898 320010 291134
rect 320246 290898 320288 291134
rect 319968 290866 320288 290898
rect 304608 273454 304928 273486
rect 304608 273218 304650 273454
rect 304886 273218 304928 273454
rect 304608 273134 304928 273218
rect 304608 272898 304650 273134
rect 304886 272898 304928 273134
rect 304608 272866 304928 272898
rect 335328 273454 335648 273486
rect 335328 273218 335370 273454
rect 335606 273218 335648 273454
rect 335328 273134 335648 273218
rect 335328 272898 335370 273134
rect 335606 272898 335648 273134
rect 335328 272866 335648 272898
rect 289248 255454 289568 255486
rect 289248 255218 289290 255454
rect 289526 255218 289568 255454
rect 289248 255134 289568 255218
rect 289248 254898 289290 255134
rect 289526 254898 289568 255134
rect 289248 254866 289568 254898
rect 319968 255454 320288 255486
rect 319968 255218 320010 255454
rect 320246 255218 320288 255454
rect 319968 255134 320288 255218
rect 319968 254898 320010 255134
rect 320246 254898 320288 255134
rect 319968 254866 320288 254898
rect 304608 237454 304928 237486
rect 304608 237218 304650 237454
rect 304886 237218 304928 237454
rect 304608 237134 304928 237218
rect 304608 236898 304650 237134
rect 304886 236898 304928 237134
rect 304608 236866 304928 236898
rect 335328 237454 335648 237486
rect 335328 237218 335370 237454
rect 335606 237218 335648 237454
rect 335328 237134 335648 237218
rect 335328 236898 335370 237134
rect 335606 236898 335648 237134
rect 335328 236866 335648 236898
rect 289248 219454 289568 219486
rect 289248 219218 289290 219454
rect 289526 219218 289568 219454
rect 289248 219134 289568 219218
rect 289248 218898 289290 219134
rect 289526 218898 289568 219134
rect 289248 218866 289568 218898
rect 319968 219454 320288 219486
rect 319968 219218 320010 219454
rect 320246 219218 320288 219454
rect 319968 219134 320288 219218
rect 319968 218898 320010 219134
rect 320246 218898 320288 219134
rect 319968 218866 320288 218898
rect 304608 201454 304928 201486
rect 304608 201218 304650 201454
rect 304886 201218 304928 201454
rect 304608 201134 304928 201218
rect 304608 200898 304650 201134
rect 304886 200898 304928 201134
rect 304608 200866 304928 200898
rect 335328 201454 335648 201486
rect 335328 201218 335370 201454
rect 335606 201218 335648 201454
rect 335328 201134 335648 201218
rect 335328 200898 335370 201134
rect 335606 200898 335648 201134
rect 335328 200866 335648 200898
rect 289248 183454 289568 183486
rect 289248 183218 289290 183454
rect 289526 183218 289568 183454
rect 289248 183134 289568 183218
rect 289248 182898 289290 183134
rect 289526 182898 289568 183134
rect 289248 182866 289568 182898
rect 319968 183454 320288 183486
rect 319968 183218 320010 183454
rect 320246 183218 320288 183454
rect 319968 183134 320288 183218
rect 319968 182898 320010 183134
rect 320246 182898 320288 183134
rect 319968 182866 320288 182898
rect 304608 165454 304928 165486
rect 304608 165218 304650 165454
rect 304886 165218 304928 165454
rect 304608 165134 304928 165218
rect 304608 164898 304650 165134
rect 304886 164898 304928 165134
rect 304608 164866 304928 164898
rect 335328 165454 335648 165486
rect 335328 165218 335370 165454
rect 335606 165218 335648 165454
rect 335328 165134 335648 165218
rect 335328 164898 335370 165134
rect 335606 164898 335648 165134
rect 335328 164866 335648 164898
rect 289248 147454 289568 147486
rect 289248 147218 289290 147454
rect 289526 147218 289568 147454
rect 289248 147134 289568 147218
rect 289248 146898 289290 147134
rect 289526 146898 289568 147134
rect 289248 146866 289568 146898
rect 319968 147454 320288 147486
rect 319968 147218 320010 147454
rect 320246 147218 320288 147454
rect 319968 147134 320288 147218
rect 319968 146898 320010 147134
rect 320246 146898 320288 147134
rect 319968 146866 320288 146898
rect 304608 129454 304928 129486
rect 304608 129218 304650 129454
rect 304886 129218 304928 129454
rect 304608 129134 304928 129218
rect 304608 128898 304650 129134
rect 304886 128898 304928 129134
rect 304608 128866 304928 128898
rect 335328 129454 335648 129486
rect 335328 129218 335370 129454
rect 335606 129218 335648 129454
rect 335328 129134 335648 129218
rect 335328 128898 335370 129134
rect 335606 128898 335648 129134
rect 335328 128866 335648 128898
rect 289248 111454 289568 111486
rect 289248 111218 289290 111454
rect 289526 111218 289568 111454
rect 289248 111134 289568 111218
rect 289248 110898 289290 111134
rect 289526 110898 289568 111134
rect 289248 110866 289568 110898
rect 319968 111454 320288 111486
rect 319968 111218 320010 111454
rect 320246 111218 320288 111454
rect 319968 111134 320288 111218
rect 319968 110898 320010 111134
rect 320246 110898 320288 111134
rect 319968 110866 320288 110898
rect 304608 93454 304928 93486
rect 304608 93218 304650 93454
rect 304886 93218 304928 93454
rect 304608 93134 304928 93218
rect 304608 92898 304650 93134
rect 304886 92898 304928 93134
rect 304608 92866 304928 92898
rect 335328 93454 335648 93486
rect 335328 93218 335370 93454
rect 335606 93218 335648 93454
rect 335328 93134 335648 93218
rect 335328 92898 335370 93134
rect 335606 92898 335648 93134
rect 335328 92866 335648 92898
rect 289248 75454 289568 75486
rect 289248 75218 289290 75454
rect 289526 75218 289568 75454
rect 289248 75134 289568 75218
rect 289248 74898 289290 75134
rect 289526 74898 289568 75134
rect 289248 74866 289568 74898
rect 319968 75454 320288 75486
rect 319968 75218 320010 75454
rect 320246 75218 320288 75454
rect 319968 75134 320288 75218
rect 319968 74898 320010 75134
rect 320246 74898 320288 75134
rect 319968 74866 320288 74898
rect 282954 32614 283574 66000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 281579 6084 281645 6085
rect 281579 6020 281580 6084
rect 281644 6020 281645 6084
rect 281579 6019 281645 6020
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 66000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 66000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 66000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 66000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 66000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 66000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 66000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 66000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 66000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 66000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 66000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 66000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 66000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 345062 6765 345122 567291
rect 346902 6901 346962 570827
rect 347514 570000 348134 600618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 348371 570756 348437 570757
rect 348371 570692 348372 570756
rect 348436 570692 348437 570756
rect 348371 570691 348437 570692
rect 347514 61174 348134 66000
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 346899 6900 346965 6901
rect 346899 6836 346900 6900
rect 346964 6836 346965 6900
rect 346899 6835 346965 6836
rect 345059 6764 345125 6765
rect 345059 6700 345060 6764
rect 345124 6700 345125 6764
rect 345059 6699 345125 6700
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 -3226 348134 24618
rect 348374 4997 348434 570691
rect 351234 570000 351854 604338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 570000 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 570000 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 570000 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 570000 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 570000 373574 590058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 570000 380414 596898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 570000 384134 600618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 570000 387854 604338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 570000 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 570000 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 570000 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 403571 570212 403637 570213
rect 403571 570148 403572 570212
rect 403636 570148 403637 570212
rect 403571 570147 403637 570148
rect 386459 567356 386525 567357
rect 386459 567292 386460 567356
rect 386524 567292 386525 567356
rect 386459 567291 386525 567292
rect 366048 561454 366368 561486
rect 366048 561218 366090 561454
rect 366326 561218 366368 561454
rect 366048 561134 366368 561218
rect 366048 560898 366090 561134
rect 366326 560898 366368 561134
rect 366048 560866 366368 560898
rect 350688 543454 351008 543486
rect 350688 543218 350730 543454
rect 350966 543218 351008 543454
rect 350688 543134 351008 543218
rect 350688 542898 350730 543134
rect 350966 542898 351008 543134
rect 350688 542866 351008 542898
rect 381408 543454 381728 543486
rect 381408 543218 381450 543454
rect 381686 543218 381728 543454
rect 381408 543134 381728 543218
rect 381408 542898 381450 543134
rect 381686 542898 381728 543134
rect 381408 542866 381728 542898
rect 366048 525454 366368 525486
rect 366048 525218 366090 525454
rect 366326 525218 366368 525454
rect 366048 525134 366368 525218
rect 366048 524898 366090 525134
rect 366326 524898 366368 525134
rect 366048 524866 366368 524898
rect 350688 507454 351008 507486
rect 350688 507218 350730 507454
rect 350966 507218 351008 507454
rect 350688 507134 351008 507218
rect 350688 506898 350730 507134
rect 350966 506898 351008 507134
rect 350688 506866 351008 506898
rect 381408 507454 381728 507486
rect 381408 507218 381450 507454
rect 381686 507218 381728 507454
rect 381408 507134 381728 507218
rect 381408 506898 381450 507134
rect 381686 506898 381728 507134
rect 381408 506866 381728 506898
rect 366048 489454 366368 489486
rect 366048 489218 366090 489454
rect 366326 489218 366368 489454
rect 366048 489134 366368 489218
rect 366048 488898 366090 489134
rect 366326 488898 366368 489134
rect 366048 488866 366368 488898
rect 350688 471454 351008 471486
rect 350688 471218 350730 471454
rect 350966 471218 351008 471454
rect 350688 471134 351008 471218
rect 350688 470898 350730 471134
rect 350966 470898 351008 471134
rect 350688 470866 351008 470898
rect 381408 471454 381728 471486
rect 381408 471218 381450 471454
rect 381686 471218 381728 471454
rect 381408 471134 381728 471218
rect 381408 470898 381450 471134
rect 381686 470898 381728 471134
rect 381408 470866 381728 470898
rect 366048 453454 366368 453486
rect 366048 453218 366090 453454
rect 366326 453218 366368 453454
rect 366048 453134 366368 453218
rect 366048 452898 366090 453134
rect 366326 452898 366368 453134
rect 366048 452866 366368 452898
rect 350688 435454 351008 435486
rect 350688 435218 350730 435454
rect 350966 435218 351008 435454
rect 350688 435134 351008 435218
rect 350688 434898 350730 435134
rect 350966 434898 351008 435134
rect 350688 434866 351008 434898
rect 381408 435454 381728 435486
rect 381408 435218 381450 435454
rect 381686 435218 381728 435454
rect 381408 435134 381728 435218
rect 381408 434898 381450 435134
rect 381686 434898 381728 435134
rect 381408 434866 381728 434898
rect 366048 417454 366368 417486
rect 366048 417218 366090 417454
rect 366326 417218 366368 417454
rect 366048 417134 366368 417218
rect 366048 416898 366090 417134
rect 366326 416898 366368 417134
rect 366048 416866 366368 416898
rect 350688 399454 351008 399486
rect 350688 399218 350730 399454
rect 350966 399218 351008 399454
rect 350688 399134 351008 399218
rect 350688 398898 350730 399134
rect 350966 398898 351008 399134
rect 350688 398866 351008 398898
rect 381408 399454 381728 399486
rect 381408 399218 381450 399454
rect 381686 399218 381728 399454
rect 381408 399134 381728 399218
rect 381408 398898 381450 399134
rect 381686 398898 381728 399134
rect 381408 398866 381728 398898
rect 366048 381454 366368 381486
rect 366048 381218 366090 381454
rect 366326 381218 366368 381454
rect 366048 381134 366368 381218
rect 366048 380898 366090 381134
rect 366326 380898 366368 381134
rect 366048 380866 366368 380898
rect 350688 363454 351008 363486
rect 350688 363218 350730 363454
rect 350966 363218 351008 363454
rect 350688 363134 351008 363218
rect 350688 362898 350730 363134
rect 350966 362898 351008 363134
rect 350688 362866 351008 362898
rect 381408 363454 381728 363486
rect 381408 363218 381450 363454
rect 381686 363218 381728 363454
rect 381408 363134 381728 363218
rect 381408 362898 381450 363134
rect 381686 362898 381728 363134
rect 381408 362866 381728 362898
rect 366048 345454 366368 345486
rect 366048 345218 366090 345454
rect 366326 345218 366368 345454
rect 366048 345134 366368 345218
rect 366048 344898 366090 345134
rect 366326 344898 366368 345134
rect 366048 344866 366368 344898
rect 350688 327454 351008 327486
rect 350688 327218 350730 327454
rect 350966 327218 351008 327454
rect 350688 327134 351008 327218
rect 350688 326898 350730 327134
rect 350966 326898 351008 327134
rect 350688 326866 351008 326898
rect 381408 327454 381728 327486
rect 381408 327218 381450 327454
rect 381686 327218 381728 327454
rect 381408 327134 381728 327218
rect 381408 326898 381450 327134
rect 381686 326898 381728 327134
rect 381408 326866 381728 326898
rect 366048 309454 366368 309486
rect 366048 309218 366090 309454
rect 366326 309218 366368 309454
rect 366048 309134 366368 309218
rect 366048 308898 366090 309134
rect 366326 308898 366368 309134
rect 366048 308866 366368 308898
rect 350688 291454 351008 291486
rect 350688 291218 350730 291454
rect 350966 291218 351008 291454
rect 350688 291134 351008 291218
rect 350688 290898 350730 291134
rect 350966 290898 351008 291134
rect 350688 290866 351008 290898
rect 381408 291454 381728 291486
rect 381408 291218 381450 291454
rect 381686 291218 381728 291454
rect 381408 291134 381728 291218
rect 381408 290898 381450 291134
rect 381686 290898 381728 291134
rect 381408 290866 381728 290898
rect 366048 273454 366368 273486
rect 366048 273218 366090 273454
rect 366326 273218 366368 273454
rect 366048 273134 366368 273218
rect 366048 272898 366090 273134
rect 366326 272898 366368 273134
rect 366048 272866 366368 272898
rect 350688 255454 351008 255486
rect 350688 255218 350730 255454
rect 350966 255218 351008 255454
rect 350688 255134 351008 255218
rect 350688 254898 350730 255134
rect 350966 254898 351008 255134
rect 350688 254866 351008 254898
rect 381408 255454 381728 255486
rect 381408 255218 381450 255454
rect 381686 255218 381728 255454
rect 381408 255134 381728 255218
rect 381408 254898 381450 255134
rect 381686 254898 381728 255134
rect 381408 254866 381728 254898
rect 366048 237454 366368 237486
rect 366048 237218 366090 237454
rect 366326 237218 366368 237454
rect 366048 237134 366368 237218
rect 366048 236898 366090 237134
rect 366326 236898 366368 237134
rect 366048 236866 366368 236898
rect 350688 219454 351008 219486
rect 350688 219218 350730 219454
rect 350966 219218 351008 219454
rect 350688 219134 351008 219218
rect 350688 218898 350730 219134
rect 350966 218898 351008 219134
rect 350688 218866 351008 218898
rect 381408 219454 381728 219486
rect 381408 219218 381450 219454
rect 381686 219218 381728 219454
rect 381408 219134 381728 219218
rect 381408 218898 381450 219134
rect 381686 218898 381728 219134
rect 381408 218866 381728 218898
rect 366048 201454 366368 201486
rect 366048 201218 366090 201454
rect 366326 201218 366368 201454
rect 366048 201134 366368 201218
rect 366048 200898 366090 201134
rect 366326 200898 366368 201134
rect 366048 200866 366368 200898
rect 350688 183454 351008 183486
rect 350688 183218 350730 183454
rect 350966 183218 351008 183454
rect 350688 183134 351008 183218
rect 350688 182898 350730 183134
rect 350966 182898 351008 183134
rect 350688 182866 351008 182898
rect 381408 183454 381728 183486
rect 381408 183218 381450 183454
rect 381686 183218 381728 183454
rect 381408 183134 381728 183218
rect 381408 182898 381450 183134
rect 381686 182898 381728 183134
rect 381408 182866 381728 182898
rect 366048 165454 366368 165486
rect 366048 165218 366090 165454
rect 366326 165218 366368 165454
rect 366048 165134 366368 165218
rect 366048 164898 366090 165134
rect 366326 164898 366368 165134
rect 366048 164866 366368 164898
rect 350688 147454 351008 147486
rect 350688 147218 350730 147454
rect 350966 147218 351008 147454
rect 350688 147134 351008 147218
rect 350688 146898 350730 147134
rect 350966 146898 351008 147134
rect 350688 146866 351008 146898
rect 381408 147454 381728 147486
rect 381408 147218 381450 147454
rect 381686 147218 381728 147454
rect 381408 147134 381728 147218
rect 381408 146898 381450 147134
rect 381686 146898 381728 147134
rect 381408 146866 381728 146898
rect 366048 129454 366368 129486
rect 366048 129218 366090 129454
rect 366326 129218 366368 129454
rect 366048 129134 366368 129218
rect 366048 128898 366090 129134
rect 366326 128898 366368 129134
rect 366048 128866 366368 128898
rect 350688 111454 351008 111486
rect 350688 111218 350730 111454
rect 350966 111218 351008 111454
rect 350688 111134 351008 111218
rect 350688 110898 350730 111134
rect 350966 110898 351008 111134
rect 350688 110866 351008 110898
rect 381408 111454 381728 111486
rect 381408 111218 381450 111454
rect 381686 111218 381728 111454
rect 381408 111134 381728 111218
rect 381408 110898 381450 111134
rect 381686 110898 381728 111134
rect 381408 110866 381728 110898
rect 366048 93454 366368 93486
rect 366048 93218 366090 93454
rect 366326 93218 366368 93454
rect 366048 93134 366368 93218
rect 366048 92898 366090 93134
rect 366326 92898 366368 93134
rect 366048 92866 366368 92898
rect 350688 75454 351008 75486
rect 350688 75218 350730 75454
rect 350966 75218 351008 75454
rect 350688 75134 351008 75218
rect 350688 74898 350730 75134
rect 350966 74898 351008 75134
rect 350688 74866 351008 74898
rect 381408 75454 381728 75486
rect 381408 75218 381450 75454
rect 381686 75218 381728 75454
rect 381408 75134 381728 75218
rect 381408 74898 381450 75134
rect 381686 74898 381728 75134
rect 381408 74866 381728 74898
rect 351234 64894 351854 66000
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 348371 4996 348437 4997
rect 348371 4932 348372 4996
rect 348436 4932 348437 4996
rect 348371 4931 348437 4932
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 66000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 66000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 66000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 66000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 66000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 66000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 61174 384134 66000
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 386462 3501 386522 567291
rect 396768 561454 397088 561486
rect 396768 561218 396810 561454
rect 397046 561218 397088 561454
rect 396768 561134 397088 561218
rect 396768 560898 396810 561134
rect 397046 560898 397088 561134
rect 396768 560866 397088 560898
rect 396768 525454 397088 525486
rect 396768 525218 396810 525454
rect 397046 525218 397088 525454
rect 396768 525134 397088 525218
rect 396768 524898 396810 525134
rect 397046 524898 397088 525134
rect 396768 524866 397088 524898
rect 396768 489454 397088 489486
rect 396768 489218 396810 489454
rect 397046 489218 397088 489454
rect 396768 489134 397088 489218
rect 396768 488898 396810 489134
rect 397046 488898 397088 489134
rect 396768 488866 397088 488898
rect 396768 453454 397088 453486
rect 396768 453218 396810 453454
rect 397046 453218 397088 453454
rect 396768 453134 397088 453218
rect 396768 452898 396810 453134
rect 397046 452898 397088 453134
rect 396768 452866 397088 452898
rect 396768 417454 397088 417486
rect 396768 417218 396810 417454
rect 397046 417218 397088 417454
rect 396768 417134 397088 417218
rect 396768 416898 396810 417134
rect 397046 416898 397088 417134
rect 396768 416866 397088 416898
rect 396768 381454 397088 381486
rect 396768 381218 396810 381454
rect 397046 381218 397088 381454
rect 396768 381134 397088 381218
rect 396768 380898 396810 381134
rect 397046 380898 397088 381134
rect 396768 380866 397088 380898
rect 396768 345454 397088 345486
rect 396768 345218 396810 345454
rect 397046 345218 397088 345454
rect 396768 345134 397088 345218
rect 396768 344898 396810 345134
rect 397046 344898 397088 345134
rect 396768 344866 397088 344898
rect 396768 309454 397088 309486
rect 396768 309218 396810 309454
rect 397046 309218 397088 309454
rect 396768 309134 397088 309218
rect 396768 308898 396810 309134
rect 397046 308898 397088 309134
rect 396768 308866 397088 308898
rect 396768 273454 397088 273486
rect 396768 273218 396810 273454
rect 397046 273218 397088 273454
rect 396768 273134 397088 273218
rect 396768 272898 396810 273134
rect 397046 272898 397088 273134
rect 396768 272866 397088 272898
rect 396768 237454 397088 237486
rect 396768 237218 396810 237454
rect 397046 237218 397088 237454
rect 396768 237134 397088 237218
rect 396768 236898 396810 237134
rect 397046 236898 397088 237134
rect 396768 236866 397088 236898
rect 396768 201454 397088 201486
rect 396768 201218 396810 201454
rect 397046 201218 397088 201454
rect 396768 201134 397088 201218
rect 396768 200898 396810 201134
rect 397046 200898 397088 201134
rect 396768 200866 397088 200898
rect 396768 165454 397088 165486
rect 396768 165218 396810 165454
rect 397046 165218 397088 165454
rect 396768 165134 397088 165218
rect 396768 164898 396810 165134
rect 397046 164898 397088 165134
rect 396768 164866 397088 164898
rect 396768 129454 397088 129486
rect 396768 129218 396810 129454
rect 397046 129218 397088 129454
rect 396768 129134 397088 129218
rect 396768 128898 396810 129134
rect 397046 128898 397088 129134
rect 396768 128866 397088 128898
rect 396768 93454 397088 93486
rect 396768 93218 396810 93454
rect 397046 93218 397088 93454
rect 396768 93134 397088 93218
rect 396768 92898 396810 93134
rect 397046 92898 397088 93134
rect 396768 92866 397088 92898
rect 387234 64894 387854 66000
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 386459 3500 386525 3501
rect 386459 3436 386460 3500
rect 386524 3436 386525 3500
rect 386459 3435 386525 3436
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 66000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 66000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 66000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 403574 6629 403634 570147
rect 405234 570000 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 570000 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 570000 416414 596898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 570000 420134 600618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 570000 423854 604338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 429147 699820 429213 699821
rect 429147 699756 429148 699820
rect 429212 699756 429213 699820
rect 429147 699755 429213 699756
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 570000 427574 572058
rect 427488 561454 427808 561486
rect 427488 561218 427530 561454
rect 427766 561218 427808 561454
rect 427488 561134 427808 561218
rect 427488 560898 427530 561134
rect 427766 560898 427808 561134
rect 427488 560866 427808 560898
rect 412128 543454 412448 543486
rect 412128 543218 412170 543454
rect 412406 543218 412448 543454
rect 412128 543134 412448 543218
rect 412128 542898 412170 543134
rect 412406 542898 412448 543134
rect 412128 542866 412448 542898
rect 427488 525454 427808 525486
rect 427488 525218 427530 525454
rect 427766 525218 427808 525454
rect 427488 525134 427808 525218
rect 427488 524898 427530 525134
rect 427766 524898 427808 525134
rect 427488 524866 427808 524898
rect 412128 507454 412448 507486
rect 412128 507218 412170 507454
rect 412406 507218 412448 507454
rect 412128 507134 412448 507218
rect 412128 506898 412170 507134
rect 412406 506898 412448 507134
rect 412128 506866 412448 506898
rect 427488 489454 427808 489486
rect 427488 489218 427530 489454
rect 427766 489218 427808 489454
rect 427488 489134 427808 489218
rect 427488 488898 427530 489134
rect 427766 488898 427808 489134
rect 427488 488866 427808 488898
rect 412128 471454 412448 471486
rect 412128 471218 412170 471454
rect 412406 471218 412448 471454
rect 412128 471134 412448 471218
rect 412128 470898 412170 471134
rect 412406 470898 412448 471134
rect 412128 470866 412448 470898
rect 427488 453454 427808 453486
rect 427488 453218 427530 453454
rect 427766 453218 427808 453454
rect 427488 453134 427808 453218
rect 427488 452898 427530 453134
rect 427766 452898 427808 453134
rect 427488 452866 427808 452898
rect 412128 435454 412448 435486
rect 412128 435218 412170 435454
rect 412406 435218 412448 435454
rect 412128 435134 412448 435218
rect 412128 434898 412170 435134
rect 412406 434898 412448 435134
rect 412128 434866 412448 434898
rect 427488 417454 427808 417486
rect 427488 417218 427530 417454
rect 427766 417218 427808 417454
rect 427488 417134 427808 417218
rect 427488 416898 427530 417134
rect 427766 416898 427808 417134
rect 427488 416866 427808 416898
rect 412128 399454 412448 399486
rect 412128 399218 412170 399454
rect 412406 399218 412448 399454
rect 412128 399134 412448 399218
rect 412128 398898 412170 399134
rect 412406 398898 412448 399134
rect 412128 398866 412448 398898
rect 427488 381454 427808 381486
rect 427488 381218 427530 381454
rect 427766 381218 427808 381454
rect 427488 381134 427808 381218
rect 427488 380898 427530 381134
rect 427766 380898 427808 381134
rect 427488 380866 427808 380898
rect 412128 363454 412448 363486
rect 412128 363218 412170 363454
rect 412406 363218 412448 363454
rect 412128 363134 412448 363218
rect 412128 362898 412170 363134
rect 412406 362898 412448 363134
rect 412128 362866 412448 362898
rect 427488 345454 427808 345486
rect 427488 345218 427530 345454
rect 427766 345218 427808 345454
rect 427488 345134 427808 345218
rect 427488 344898 427530 345134
rect 427766 344898 427808 345134
rect 427488 344866 427808 344898
rect 412128 327454 412448 327486
rect 412128 327218 412170 327454
rect 412406 327218 412448 327454
rect 412128 327134 412448 327218
rect 412128 326898 412170 327134
rect 412406 326898 412448 327134
rect 412128 326866 412448 326898
rect 427488 309454 427808 309486
rect 427488 309218 427530 309454
rect 427766 309218 427808 309454
rect 427488 309134 427808 309218
rect 427488 308898 427530 309134
rect 427766 308898 427808 309134
rect 427488 308866 427808 308898
rect 412128 291454 412448 291486
rect 412128 291218 412170 291454
rect 412406 291218 412448 291454
rect 412128 291134 412448 291218
rect 412128 290898 412170 291134
rect 412406 290898 412448 291134
rect 412128 290866 412448 290898
rect 427488 273454 427808 273486
rect 427488 273218 427530 273454
rect 427766 273218 427808 273454
rect 427488 273134 427808 273218
rect 427488 272898 427530 273134
rect 427766 272898 427808 273134
rect 427488 272866 427808 272898
rect 412128 255454 412448 255486
rect 412128 255218 412170 255454
rect 412406 255218 412448 255454
rect 412128 255134 412448 255218
rect 412128 254898 412170 255134
rect 412406 254898 412448 255134
rect 412128 254866 412448 254898
rect 427488 237454 427808 237486
rect 427488 237218 427530 237454
rect 427766 237218 427808 237454
rect 427488 237134 427808 237218
rect 427488 236898 427530 237134
rect 427766 236898 427808 237134
rect 427488 236866 427808 236898
rect 412128 219454 412448 219486
rect 412128 219218 412170 219454
rect 412406 219218 412448 219454
rect 412128 219134 412448 219218
rect 412128 218898 412170 219134
rect 412406 218898 412448 219134
rect 412128 218866 412448 218898
rect 427488 201454 427808 201486
rect 427488 201218 427530 201454
rect 427766 201218 427808 201454
rect 427488 201134 427808 201218
rect 427488 200898 427530 201134
rect 427766 200898 427808 201134
rect 427488 200866 427808 200898
rect 412128 183454 412448 183486
rect 412128 183218 412170 183454
rect 412406 183218 412448 183454
rect 412128 183134 412448 183218
rect 412128 182898 412170 183134
rect 412406 182898 412448 183134
rect 412128 182866 412448 182898
rect 427488 165454 427808 165486
rect 427488 165218 427530 165454
rect 427766 165218 427808 165454
rect 427488 165134 427808 165218
rect 427488 164898 427530 165134
rect 427766 164898 427808 165134
rect 427488 164866 427808 164898
rect 412128 147454 412448 147486
rect 412128 147218 412170 147454
rect 412406 147218 412448 147454
rect 412128 147134 412448 147218
rect 412128 146898 412170 147134
rect 412406 146898 412448 147134
rect 412128 146866 412448 146898
rect 427488 129454 427808 129486
rect 427488 129218 427530 129454
rect 427766 129218 427808 129454
rect 427488 129134 427808 129218
rect 427488 128898 427530 129134
rect 427766 128898 427808 129134
rect 427488 128866 427808 128898
rect 412128 111454 412448 111486
rect 412128 111218 412170 111454
rect 412406 111218 412448 111454
rect 412128 111134 412448 111218
rect 412128 110898 412170 111134
rect 412406 110898 412448 111134
rect 412128 110866 412448 110898
rect 427488 93454 427808 93486
rect 427488 93218 427530 93454
rect 427766 93218 427808 93454
rect 427488 93134 427808 93218
rect 427488 92898 427530 93134
rect 427766 92898 427808 93134
rect 427488 92866 427808 92898
rect 412128 75454 412448 75486
rect 412128 75218 412170 75454
rect 412406 75218 412448 75454
rect 412128 75134 412448 75218
rect 412128 74898 412170 75134
rect 412406 74898 412448 75134
rect 412128 74866 412448 74898
rect 429150 67557 429210 699755
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 570000 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 570000 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 570000 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 570000 445574 590058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 570000 452414 596898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 570000 456134 600618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 570000 459854 604338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 570000 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 570000 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 570000 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 570000 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 570000 481574 590058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 570000 488414 596898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 570000 492134 600618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 570000 495854 604338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 570000 499574 572058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 570000 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 570000 510134 582618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 570000 513854 586338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 570000 517574 590058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 570000 524414 596898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 570000 528134 600618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 570000 531854 604338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 570000 535574 572058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 570000 542414 578898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 570000 546134 582618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 570000 549854 586338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 570000 553574 590058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 570000 560414 596898
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 570000 564134 600618
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 570000 567854 604338
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 570000 571574 572058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 440187 567356 440253 567357
rect 440187 567292 440188 567356
rect 440252 567292 440253 567356
rect 440187 567291 440253 567292
rect 460979 567356 461045 567357
rect 460979 567292 460980 567356
rect 461044 567292 461045 567356
rect 460979 567291 461045 567292
rect 481771 567356 481837 567357
rect 481771 567292 481772 567356
rect 481836 567292 481837 567356
rect 481771 567291 481837 567292
rect 539547 567356 539613 567357
rect 539547 567292 539548 567356
rect 539612 567292 539613 567356
rect 539547 567291 539613 567292
rect 550771 567356 550837 567357
rect 550771 567292 550772 567356
rect 550836 567292 550837 567356
rect 550771 567291 550837 567292
rect 429147 67556 429213 67557
rect 429147 67492 429148 67556
rect 429212 67492 429213 67556
rect 429147 67491 429213 67492
rect 405234 46894 405854 66000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 401514 -2266 402134 6618
rect 403571 6628 403637 6629
rect 403571 6564 403572 6628
rect 403636 6564 403637 6628
rect 403571 6563 403637 6564
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 66000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 66000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 61174 420134 66000
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 64894 423854 66000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 66000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 66000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 66000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 440190 6357 440250 567291
rect 458208 561454 458528 561486
rect 458208 561218 458250 561454
rect 458486 561218 458528 561454
rect 458208 561134 458528 561218
rect 458208 560898 458250 561134
rect 458486 560898 458528 561134
rect 458208 560866 458528 560898
rect 442848 543454 443168 543486
rect 442848 543218 442890 543454
rect 443126 543218 443168 543454
rect 442848 543134 443168 543218
rect 442848 542898 442890 543134
rect 443126 542898 443168 543134
rect 442848 542866 443168 542898
rect 458208 525454 458528 525486
rect 458208 525218 458250 525454
rect 458486 525218 458528 525454
rect 458208 525134 458528 525218
rect 458208 524898 458250 525134
rect 458486 524898 458528 525134
rect 458208 524866 458528 524898
rect 442848 507454 443168 507486
rect 442848 507218 442890 507454
rect 443126 507218 443168 507454
rect 442848 507134 443168 507218
rect 442848 506898 442890 507134
rect 443126 506898 443168 507134
rect 442848 506866 443168 506898
rect 458208 489454 458528 489486
rect 458208 489218 458250 489454
rect 458486 489218 458528 489454
rect 458208 489134 458528 489218
rect 458208 488898 458250 489134
rect 458486 488898 458528 489134
rect 458208 488866 458528 488898
rect 442848 471454 443168 471486
rect 442848 471218 442890 471454
rect 443126 471218 443168 471454
rect 442848 471134 443168 471218
rect 442848 470898 442890 471134
rect 443126 470898 443168 471134
rect 442848 470866 443168 470898
rect 458208 453454 458528 453486
rect 458208 453218 458250 453454
rect 458486 453218 458528 453454
rect 458208 453134 458528 453218
rect 458208 452898 458250 453134
rect 458486 452898 458528 453134
rect 458208 452866 458528 452898
rect 442848 435454 443168 435486
rect 442848 435218 442890 435454
rect 443126 435218 443168 435454
rect 442848 435134 443168 435218
rect 442848 434898 442890 435134
rect 443126 434898 443168 435134
rect 442848 434866 443168 434898
rect 458208 417454 458528 417486
rect 458208 417218 458250 417454
rect 458486 417218 458528 417454
rect 458208 417134 458528 417218
rect 458208 416898 458250 417134
rect 458486 416898 458528 417134
rect 458208 416866 458528 416898
rect 442848 399454 443168 399486
rect 442848 399218 442890 399454
rect 443126 399218 443168 399454
rect 442848 399134 443168 399218
rect 442848 398898 442890 399134
rect 443126 398898 443168 399134
rect 442848 398866 443168 398898
rect 458208 381454 458528 381486
rect 458208 381218 458250 381454
rect 458486 381218 458528 381454
rect 458208 381134 458528 381218
rect 458208 380898 458250 381134
rect 458486 380898 458528 381134
rect 458208 380866 458528 380898
rect 442848 363454 443168 363486
rect 442848 363218 442890 363454
rect 443126 363218 443168 363454
rect 442848 363134 443168 363218
rect 442848 362898 442890 363134
rect 443126 362898 443168 363134
rect 442848 362866 443168 362898
rect 458208 345454 458528 345486
rect 458208 345218 458250 345454
rect 458486 345218 458528 345454
rect 458208 345134 458528 345218
rect 458208 344898 458250 345134
rect 458486 344898 458528 345134
rect 458208 344866 458528 344898
rect 442848 327454 443168 327486
rect 442848 327218 442890 327454
rect 443126 327218 443168 327454
rect 442848 327134 443168 327218
rect 442848 326898 442890 327134
rect 443126 326898 443168 327134
rect 442848 326866 443168 326898
rect 458208 309454 458528 309486
rect 458208 309218 458250 309454
rect 458486 309218 458528 309454
rect 458208 309134 458528 309218
rect 458208 308898 458250 309134
rect 458486 308898 458528 309134
rect 458208 308866 458528 308898
rect 442848 291454 443168 291486
rect 442848 291218 442890 291454
rect 443126 291218 443168 291454
rect 442848 291134 443168 291218
rect 442848 290898 442890 291134
rect 443126 290898 443168 291134
rect 442848 290866 443168 290898
rect 458208 273454 458528 273486
rect 458208 273218 458250 273454
rect 458486 273218 458528 273454
rect 458208 273134 458528 273218
rect 458208 272898 458250 273134
rect 458486 272898 458528 273134
rect 458208 272866 458528 272898
rect 442848 255454 443168 255486
rect 442848 255218 442890 255454
rect 443126 255218 443168 255454
rect 442848 255134 443168 255218
rect 442848 254898 442890 255134
rect 443126 254898 443168 255134
rect 442848 254866 443168 254898
rect 458208 237454 458528 237486
rect 458208 237218 458250 237454
rect 458486 237218 458528 237454
rect 458208 237134 458528 237218
rect 458208 236898 458250 237134
rect 458486 236898 458528 237134
rect 458208 236866 458528 236898
rect 442848 219454 443168 219486
rect 442848 219218 442890 219454
rect 443126 219218 443168 219454
rect 442848 219134 443168 219218
rect 442848 218898 442890 219134
rect 443126 218898 443168 219134
rect 442848 218866 443168 218898
rect 458208 201454 458528 201486
rect 458208 201218 458250 201454
rect 458486 201218 458528 201454
rect 458208 201134 458528 201218
rect 458208 200898 458250 201134
rect 458486 200898 458528 201134
rect 458208 200866 458528 200898
rect 442848 183454 443168 183486
rect 442848 183218 442890 183454
rect 443126 183218 443168 183454
rect 442848 183134 443168 183218
rect 442848 182898 442890 183134
rect 443126 182898 443168 183134
rect 442848 182866 443168 182898
rect 458208 165454 458528 165486
rect 458208 165218 458250 165454
rect 458486 165218 458528 165454
rect 458208 165134 458528 165218
rect 458208 164898 458250 165134
rect 458486 164898 458528 165134
rect 458208 164866 458528 164898
rect 442848 147454 443168 147486
rect 442848 147218 442890 147454
rect 443126 147218 443168 147454
rect 442848 147134 443168 147218
rect 442848 146898 442890 147134
rect 443126 146898 443168 147134
rect 442848 146866 443168 146898
rect 458208 129454 458528 129486
rect 458208 129218 458250 129454
rect 458486 129218 458528 129454
rect 458208 129134 458528 129218
rect 458208 128898 458250 129134
rect 458486 128898 458528 129134
rect 458208 128866 458528 128898
rect 442848 111454 443168 111486
rect 442848 111218 442890 111454
rect 443126 111218 443168 111454
rect 442848 111134 443168 111218
rect 442848 110898 442890 111134
rect 443126 110898 443168 111134
rect 442848 110866 443168 110898
rect 458208 93454 458528 93486
rect 458208 93218 458250 93454
rect 458486 93218 458528 93454
rect 458208 93134 458528 93218
rect 458208 92898 458250 93134
rect 458486 92898 458528 93134
rect 458208 92866 458528 92898
rect 442848 75454 443168 75486
rect 442848 75218 442890 75454
rect 443126 75218 443168 75454
rect 442848 75134 443168 75218
rect 442848 74898 442890 75134
rect 443126 74898 443168 75134
rect 442848 74866 443168 74898
rect 441234 46894 441854 66000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 440187 6356 440253 6357
rect 440187 6292 440188 6356
rect 440252 6292 440253 6356
rect 440187 6291 440253 6292
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 66000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 66000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 61174 456134 66000
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 64894 459854 66000
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 460982 6493 461042 567291
rect 473568 543454 473888 543486
rect 473568 543218 473610 543454
rect 473846 543218 473888 543454
rect 473568 543134 473888 543218
rect 473568 542898 473610 543134
rect 473846 542898 473888 543134
rect 473568 542866 473888 542898
rect 473568 507454 473888 507486
rect 473568 507218 473610 507454
rect 473846 507218 473888 507454
rect 473568 507134 473888 507218
rect 473568 506898 473610 507134
rect 473846 506898 473888 507134
rect 473568 506866 473888 506898
rect 473568 471454 473888 471486
rect 473568 471218 473610 471454
rect 473846 471218 473888 471454
rect 473568 471134 473888 471218
rect 473568 470898 473610 471134
rect 473846 470898 473888 471134
rect 473568 470866 473888 470898
rect 473568 435454 473888 435486
rect 473568 435218 473610 435454
rect 473846 435218 473888 435454
rect 473568 435134 473888 435218
rect 473568 434898 473610 435134
rect 473846 434898 473888 435134
rect 473568 434866 473888 434898
rect 473568 399454 473888 399486
rect 473568 399218 473610 399454
rect 473846 399218 473888 399454
rect 473568 399134 473888 399218
rect 473568 398898 473610 399134
rect 473846 398898 473888 399134
rect 473568 398866 473888 398898
rect 473568 363454 473888 363486
rect 473568 363218 473610 363454
rect 473846 363218 473888 363454
rect 473568 363134 473888 363218
rect 473568 362898 473610 363134
rect 473846 362898 473888 363134
rect 473568 362866 473888 362898
rect 473568 327454 473888 327486
rect 473568 327218 473610 327454
rect 473846 327218 473888 327454
rect 473568 327134 473888 327218
rect 473568 326898 473610 327134
rect 473846 326898 473888 327134
rect 473568 326866 473888 326898
rect 473568 291454 473888 291486
rect 473568 291218 473610 291454
rect 473846 291218 473888 291454
rect 473568 291134 473888 291218
rect 473568 290898 473610 291134
rect 473846 290898 473888 291134
rect 473568 290866 473888 290898
rect 473568 255454 473888 255486
rect 473568 255218 473610 255454
rect 473846 255218 473888 255454
rect 473568 255134 473888 255218
rect 473568 254898 473610 255134
rect 473846 254898 473888 255134
rect 473568 254866 473888 254898
rect 473568 219454 473888 219486
rect 473568 219218 473610 219454
rect 473846 219218 473888 219454
rect 473568 219134 473888 219218
rect 473568 218898 473610 219134
rect 473846 218898 473888 219134
rect 473568 218866 473888 218898
rect 473568 183454 473888 183486
rect 473568 183218 473610 183454
rect 473846 183218 473888 183454
rect 473568 183134 473888 183218
rect 473568 182898 473610 183134
rect 473846 182898 473888 183134
rect 473568 182866 473888 182898
rect 473568 147454 473888 147486
rect 473568 147218 473610 147454
rect 473846 147218 473888 147454
rect 473568 147134 473888 147218
rect 473568 146898 473610 147134
rect 473846 146898 473888 147134
rect 473568 146866 473888 146898
rect 473568 111454 473888 111486
rect 473568 111218 473610 111454
rect 473846 111218 473888 111454
rect 473568 111134 473888 111218
rect 473568 110898 473610 111134
rect 473846 110898 473888 111134
rect 473568 110866 473888 110898
rect 473568 75454 473888 75486
rect 473568 75218 473610 75454
rect 473846 75218 473888 75454
rect 473568 75134 473888 75218
rect 473568 74898 473610 75134
rect 473846 74898 473888 75134
rect 473568 74866 473888 74898
rect 462954 32614 463574 66000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 460979 6492 461045 6493
rect 460979 6428 460980 6492
rect 461044 6428 461045 6492
rect 460979 6427 461045 6428
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 66000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 66000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 66000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 66000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 481774 6221 481834 567291
rect 488928 561454 489248 561486
rect 488928 561218 488970 561454
rect 489206 561218 489248 561454
rect 488928 561134 489248 561218
rect 488928 560898 488970 561134
rect 489206 560898 489248 561134
rect 488928 560866 489248 560898
rect 519648 561454 519968 561486
rect 519648 561218 519690 561454
rect 519926 561218 519968 561454
rect 519648 561134 519968 561218
rect 519648 560898 519690 561134
rect 519926 560898 519968 561134
rect 519648 560866 519968 560898
rect 504288 543454 504608 543486
rect 504288 543218 504330 543454
rect 504566 543218 504608 543454
rect 504288 543134 504608 543218
rect 504288 542898 504330 543134
rect 504566 542898 504608 543134
rect 504288 542866 504608 542898
rect 535008 543454 535328 543486
rect 535008 543218 535050 543454
rect 535286 543218 535328 543454
rect 535008 543134 535328 543218
rect 535008 542898 535050 543134
rect 535286 542898 535328 543134
rect 535008 542866 535328 542898
rect 488928 525454 489248 525486
rect 488928 525218 488970 525454
rect 489206 525218 489248 525454
rect 488928 525134 489248 525218
rect 488928 524898 488970 525134
rect 489206 524898 489248 525134
rect 488928 524866 489248 524898
rect 519648 525454 519968 525486
rect 519648 525218 519690 525454
rect 519926 525218 519968 525454
rect 519648 525134 519968 525218
rect 519648 524898 519690 525134
rect 519926 524898 519968 525134
rect 519648 524866 519968 524898
rect 504288 507454 504608 507486
rect 504288 507218 504330 507454
rect 504566 507218 504608 507454
rect 504288 507134 504608 507218
rect 504288 506898 504330 507134
rect 504566 506898 504608 507134
rect 504288 506866 504608 506898
rect 535008 507454 535328 507486
rect 535008 507218 535050 507454
rect 535286 507218 535328 507454
rect 535008 507134 535328 507218
rect 535008 506898 535050 507134
rect 535286 506898 535328 507134
rect 535008 506866 535328 506898
rect 488928 489454 489248 489486
rect 488928 489218 488970 489454
rect 489206 489218 489248 489454
rect 488928 489134 489248 489218
rect 488928 488898 488970 489134
rect 489206 488898 489248 489134
rect 488928 488866 489248 488898
rect 519648 489454 519968 489486
rect 519648 489218 519690 489454
rect 519926 489218 519968 489454
rect 519648 489134 519968 489218
rect 519648 488898 519690 489134
rect 519926 488898 519968 489134
rect 519648 488866 519968 488898
rect 504288 471454 504608 471486
rect 504288 471218 504330 471454
rect 504566 471218 504608 471454
rect 504288 471134 504608 471218
rect 504288 470898 504330 471134
rect 504566 470898 504608 471134
rect 504288 470866 504608 470898
rect 535008 471454 535328 471486
rect 535008 471218 535050 471454
rect 535286 471218 535328 471454
rect 535008 471134 535328 471218
rect 535008 470898 535050 471134
rect 535286 470898 535328 471134
rect 535008 470866 535328 470898
rect 488928 453454 489248 453486
rect 488928 453218 488970 453454
rect 489206 453218 489248 453454
rect 488928 453134 489248 453218
rect 488928 452898 488970 453134
rect 489206 452898 489248 453134
rect 488928 452866 489248 452898
rect 519648 453454 519968 453486
rect 519648 453218 519690 453454
rect 519926 453218 519968 453454
rect 519648 453134 519968 453218
rect 519648 452898 519690 453134
rect 519926 452898 519968 453134
rect 519648 452866 519968 452898
rect 504288 435454 504608 435486
rect 504288 435218 504330 435454
rect 504566 435218 504608 435454
rect 504288 435134 504608 435218
rect 504288 434898 504330 435134
rect 504566 434898 504608 435134
rect 504288 434866 504608 434898
rect 535008 435454 535328 435486
rect 535008 435218 535050 435454
rect 535286 435218 535328 435454
rect 535008 435134 535328 435218
rect 535008 434898 535050 435134
rect 535286 434898 535328 435134
rect 535008 434866 535328 434898
rect 488928 417454 489248 417486
rect 488928 417218 488970 417454
rect 489206 417218 489248 417454
rect 488928 417134 489248 417218
rect 488928 416898 488970 417134
rect 489206 416898 489248 417134
rect 488928 416866 489248 416898
rect 519648 417454 519968 417486
rect 519648 417218 519690 417454
rect 519926 417218 519968 417454
rect 519648 417134 519968 417218
rect 519648 416898 519690 417134
rect 519926 416898 519968 417134
rect 519648 416866 519968 416898
rect 504288 399454 504608 399486
rect 504288 399218 504330 399454
rect 504566 399218 504608 399454
rect 504288 399134 504608 399218
rect 504288 398898 504330 399134
rect 504566 398898 504608 399134
rect 504288 398866 504608 398898
rect 535008 399454 535328 399486
rect 535008 399218 535050 399454
rect 535286 399218 535328 399454
rect 535008 399134 535328 399218
rect 535008 398898 535050 399134
rect 535286 398898 535328 399134
rect 535008 398866 535328 398898
rect 488928 381454 489248 381486
rect 488928 381218 488970 381454
rect 489206 381218 489248 381454
rect 488928 381134 489248 381218
rect 488928 380898 488970 381134
rect 489206 380898 489248 381134
rect 488928 380866 489248 380898
rect 519648 381454 519968 381486
rect 519648 381218 519690 381454
rect 519926 381218 519968 381454
rect 519648 381134 519968 381218
rect 519648 380898 519690 381134
rect 519926 380898 519968 381134
rect 519648 380866 519968 380898
rect 504288 363454 504608 363486
rect 504288 363218 504330 363454
rect 504566 363218 504608 363454
rect 504288 363134 504608 363218
rect 504288 362898 504330 363134
rect 504566 362898 504608 363134
rect 504288 362866 504608 362898
rect 535008 363454 535328 363486
rect 535008 363218 535050 363454
rect 535286 363218 535328 363454
rect 535008 363134 535328 363218
rect 535008 362898 535050 363134
rect 535286 362898 535328 363134
rect 535008 362866 535328 362898
rect 488928 345454 489248 345486
rect 488928 345218 488970 345454
rect 489206 345218 489248 345454
rect 488928 345134 489248 345218
rect 488928 344898 488970 345134
rect 489206 344898 489248 345134
rect 488928 344866 489248 344898
rect 519648 345454 519968 345486
rect 519648 345218 519690 345454
rect 519926 345218 519968 345454
rect 519648 345134 519968 345218
rect 519648 344898 519690 345134
rect 519926 344898 519968 345134
rect 519648 344866 519968 344898
rect 504288 327454 504608 327486
rect 504288 327218 504330 327454
rect 504566 327218 504608 327454
rect 504288 327134 504608 327218
rect 504288 326898 504330 327134
rect 504566 326898 504608 327134
rect 504288 326866 504608 326898
rect 535008 327454 535328 327486
rect 535008 327218 535050 327454
rect 535286 327218 535328 327454
rect 535008 327134 535328 327218
rect 535008 326898 535050 327134
rect 535286 326898 535328 327134
rect 535008 326866 535328 326898
rect 488928 309454 489248 309486
rect 488928 309218 488970 309454
rect 489206 309218 489248 309454
rect 488928 309134 489248 309218
rect 488928 308898 488970 309134
rect 489206 308898 489248 309134
rect 488928 308866 489248 308898
rect 519648 309454 519968 309486
rect 519648 309218 519690 309454
rect 519926 309218 519968 309454
rect 519648 309134 519968 309218
rect 519648 308898 519690 309134
rect 519926 308898 519968 309134
rect 519648 308866 519968 308898
rect 504288 291454 504608 291486
rect 504288 291218 504330 291454
rect 504566 291218 504608 291454
rect 504288 291134 504608 291218
rect 504288 290898 504330 291134
rect 504566 290898 504608 291134
rect 504288 290866 504608 290898
rect 535008 291454 535328 291486
rect 535008 291218 535050 291454
rect 535286 291218 535328 291454
rect 535008 291134 535328 291218
rect 535008 290898 535050 291134
rect 535286 290898 535328 291134
rect 535008 290866 535328 290898
rect 488928 273454 489248 273486
rect 488928 273218 488970 273454
rect 489206 273218 489248 273454
rect 488928 273134 489248 273218
rect 488928 272898 488970 273134
rect 489206 272898 489248 273134
rect 488928 272866 489248 272898
rect 519648 273454 519968 273486
rect 519648 273218 519690 273454
rect 519926 273218 519968 273454
rect 519648 273134 519968 273218
rect 519648 272898 519690 273134
rect 519926 272898 519968 273134
rect 519648 272866 519968 272898
rect 504288 255454 504608 255486
rect 504288 255218 504330 255454
rect 504566 255218 504608 255454
rect 504288 255134 504608 255218
rect 504288 254898 504330 255134
rect 504566 254898 504608 255134
rect 504288 254866 504608 254898
rect 535008 255454 535328 255486
rect 535008 255218 535050 255454
rect 535286 255218 535328 255454
rect 535008 255134 535328 255218
rect 535008 254898 535050 255134
rect 535286 254898 535328 255134
rect 535008 254866 535328 254898
rect 488928 237454 489248 237486
rect 488928 237218 488970 237454
rect 489206 237218 489248 237454
rect 488928 237134 489248 237218
rect 488928 236898 488970 237134
rect 489206 236898 489248 237134
rect 488928 236866 489248 236898
rect 519648 237454 519968 237486
rect 519648 237218 519690 237454
rect 519926 237218 519968 237454
rect 519648 237134 519968 237218
rect 519648 236898 519690 237134
rect 519926 236898 519968 237134
rect 519648 236866 519968 236898
rect 504288 219454 504608 219486
rect 504288 219218 504330 219454
rect 504566 219218 504608 219454
rect 504288 219134 504608 219218
rect 504288 218898 504330 219134
rect 504566 218898 504608 219134
rect 504288 218866 504608 218898
rect 535008 219454 535328 219486
rect 535008 219218 535050 219454
rect 535286 219218 535328 219454
rect 535008 219134 535328 219218
rect 535008 218898 535050 219134
rect 535286 218898 535328 219134
rect 535008 218866 535328 218898
rect 488928 201454 489248 201486
rect 488928 201218 488970 201454
rect 489206 201218 489248 201454
rect 488928 201134 489248 201218
rect 488928 200898 488970 201134
rect 489206 200898 489248 201134
rect 488928 200866 489248 200898
rect 519648 201454 519968 201486
rect 519648 201218 519690 201454
rect 519926 201218 519968 201454
rect 519648 201134 519968 201218
rect 519648 200898 519690 201134
rect 519926 200898 519968 201134
rect 519648 200866 519968 200898
rect 504288 183454 504608 183486
rect 504288 183218 504330 183454
rect 504566 183218 504608 183454
rect 504288 183134 504608 183218
rect 504288 182898 504330 183134
rect 504566 182898 504608 183134
rect 504288 182866 504608 182898
rect 535008 183454 535328 183486
rect 535008 183218 535050 183454
rect 535286 183218 535328 183454
rect 535008 183134 535328 183218
rect 535008 182898 535050 183134
rect 535286 182898 535328 183134
rect 535008 182866 535328 182898
rect 488928 165454 489248 165486
rect 488928 165218 488970 165454
rect 489206 165218 489248 165454
rect 488928 165134 489248 165218
rect 488928 164898 488970 165134
rect 489206 164898 489248 165134
rect 488928 164866 489248 164898
rect 519648 165454 519968 165486
rect 519648 165218 519690 165454
rect 519926 165218 519968 165454
rect 519648 165134 519968 165218
rect 519648 164898 519690 165134
rect 519926 164898 519968 165134
rect 519648 164866 519968 164898
rect 504288 147454 504608 147486
rect 504288 147218 504330 147454
rect 504566 147218 504608 147454
rect 504288 147134 504608 147218
rect 504288 146898 504330 147134
rect 504566 146898 504608 147134
rect 504288 146866 504608 146898
rect 535008 147454 535328 147486
rect 535008 147218 535050 147454
rect 535286 147218 535328 147454
rect 535008 147134 535328 147218
rect 535008 146898 535050 147134
rect 535286 146898 535328 147134
rect 535008 146866 535328 146898
rect 488928 129454 489248 129486
rect 488928 129218 488970 129454
rect 489206 129218 489248 129454
rect 488928 129134 489248 129218
rect 488928 128898 488970 129134
rect 489206 128898 489248 129134
rect 488928 128866 489248 128898
rect 519648 129454 519968 129486
rect 519648 129218 519690 129454
rect 519926 129218 519968 129454
rect 519648 129134 519968 129218
rect 519648 128898 519690 129134
rect 519926 128898 519968 129134
rect 519648 128866 519968 128898
rect 504288 111454 504608 111486
rect 504288 111218 504330 111454
rect 504566 111218 504608 111454
rect 504288 111134 504608 111218
rect 504288 110898 504330 111134
rect 504566 110898 504608 111134
rect 504288 110866 504608 110898
rect 535008 111454 535328 111486
rect 535008 111218 535050 111454
rect 535286 111218 535328 111454
rect 535008 111134 535328 111218
rect 535008 110898 535050 111134
rect 535286 110898 535328 111134
rect 535008 110866 535328 110898
rect 488928 93454 489248 93486
rect 488928 93218 488970 93454
rect 489206 93218 489248 93454
rect 488928 93134 489248 93218
rect 488928 92898 488970 93134
rect 489206 92898 489248 93134
rect 488928 92866 489248 92898
rect 519648 93454 519968 93486
rect 519648 93218 519690 93454
rect 519926 93218 519968 93454
rect 519648 93134 519968 93218
rect 519648 92898 519690 93134
rect 519926 92898 519968 93134
rect 519648 92866 519968 92898
rect 504288 75454 504608 75486
rect 504288 75218 504330 75454
rect 504566 75218 504608 75454
rect 504288 75134 504608 75218
rect 504288 74898 504330 75134
rect 504566 74898 504608 75134
rect 504288 74866 504608 74898
rect 535008 75454 535328 75486
rect 535008 75218 535050 75454
rect 535286 75218 535328 75454
rect 535008 75134 535328 75218
rect 535008 74898 535050 75134
rect 535286 74898 535328 75134
rect 535008 74866 535328 74898
rect 487794 57454 488414 66000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 481771 6220 481837 6221
rect 481771 6156 481772 6220
rect 481836 6156 481837 6220
rect 481771 6155 481837 6156
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 61174 492134 66000
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 64894 495854 66000
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 66000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 66000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 66000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 66000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 66000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 66000
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 61174 528134 66000
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 64894 531854 66000
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 66000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 539550 3365 539610 567291
rect 550368 561454 550688 561486
rect 550368 561218 550410 561454
rect 550646 561218 550688 561454
rect 550368 561134 550688 561218
rect 550368 560898 550410 561134
rect 550646 560898 550688 561134
rect 550368 560866 550688 560898
rect 550368 525454 550688 525486
rect 550368 525218 550410 525454
rect 550646 525218 550688 525454
rect 550368 525134 550688 525218
rect 550368 524898 550410 525134
rect 550646 524898 550688 525134
rect 550368 524866 550688 524898
rect 550368 489454 550688 489486
rect 550368 489218 550410 489454
rect 550646 489218 550688 489454
rect 550368 489134 550688 489218
rect 550368 488898 550410 489134
rect 550646 488898 550688 489134
rect 550368 488866 550688 488898
rect 550368 453454 550688 453486
rect 550368 453218 550410 453454
rect 550646 453218 550688 453454
rect 550368 453134 550688 453218
rect 550368 452898 550410 453134
rect 550646 452898 550688 453134
rect 550368 452866 550688 452898
rect 550368 417454 550688 417486
rect 550368 417218 550410 417454
rect 550646 417218 550688 417454
rect 550368 417134 550688 417218
rect 550368 416898 550410 417134
rect 550646 416898 550688 417134
rect 550368 416866 550688 416898
rect 550368 381454 550688 381486
rect 550368 381218 550410 381454
rect 550646 381218 550688 381454
rect 550368 381134 550688 381218
rect 550368 380898 550410 381134
rect 550646 380898 550688 381134
rect 550368 380866 550688 380898
rect 550368 345454 550688 345486
rect 550368 345218 550410 345454
rect 550646 345218 550688 345454
rect 550368 345134 550688 345218
rect 550368 344898 550410 345134
rect 550646 344898 550688 345134
rect 550368 344866 550688 344898
rect 550368 309454 550688 309486
rect 550368 309218 550410 309454
rect 550646 309218 550688 309454
rect 550368 309134 550688 309218
rect 550368 308898 550410 309134
rect 550646 308898 550688 309134
rect 550368 308866 550688 308898
rect 550368 273454 550688 273486
rect 550368 273218 550410 273454
rect 550646 273218 550688 273454
rect 550368 273134 550688 273218
rect 550368 272898 550410 273134
rect 550646 272898 550688 273134
rect 550368 272866 550688 272898
rect 550368 237454 550688 237486
rect 550368 237218 550410 237454
rect 550646 237218 550688 237454
rect 550368 237134 550688 237218
rect 550368 236898 550410 237134
rect 550646 236898 550688 237134
rect 550368 236866 550688 236898
rect 550368 201454 550688 201486
rect 550368 201218 550410 201454
rect 550646 201218 550688 201454
rect 550368 201134 550688 201218
rect 550368 200898 550410 201134
rect 550646 200898 550688 201134
rect 550368 200866 550688 200898
rect 550368 165454 550688 165486
rect 550368 165218 550410 165454
rect 550646 165218 550688 165454
rect 550368 165134 550688 165218
rect 550368 164898 550410 165134
rect 550646 164898 550688 165134
rect 550368 164866 550688 164898
rect 550368 129454 550688 129486
rect 550368 129218 550410 129454
rect 550646 129218 550688 129454
rect 550368 129134 550688 129218
rect 550368 128898 550410 129134
rect 550646 128898 550688 129134
rect 550368 128866 550688 128898
rect 550368 93454 550688 93486
rect 550368 93218 550410 93454
rect 550646 93218 550688 93454
rect 550368 93134 550688 93218
rect 550368 92898 550410 93134
rect 550646 92898 550688 93134
rect 550368 92866 550688 92898
rect 541794 39454 542414 66000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 539547 3364 539613 3365
rect 539547 3300 539548 3364
rect 539612 3300 539613 3364
rect 539547 3299 539613 3300
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 66000
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 46894 549854 66000
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 550774 4861 550834 567291
rect 565728 543454 566048 543486
rect 565728 543218 565770 543454
rect 566006 543218 566048 543454
rect 565728 543134 566048 543218
rect 565728 542898 565770 543134
rect 566006 542898 566048 543134
rect 565728 542866 566048 542898
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 565728 507454 566048 507486
rect 565728 507218 565770 507454
rect 566006 507218 566048 507454
rect 565728 507134 566048 507218
rect 565728 506898 565770 507134
rect 566006 506898 566048 507134
rect 565728 506866 566048 506898
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 565728 471454 566048 471486
rect 565728 471218 565770 471454
rect 566006 471218 566048 471454
rect 565728 471134 566048 471218
rect 565728 470898 565770 471134
rect 566006 470898 566048 471134
rect 565728 470866 566048 470898
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 565728 435454 566048 435486
rect 565728 435218 565770 435454
rect 566006 435218 566048 435454
rect 565728 435134 566048 435218
rect 565728 434898 565770 435134
rect 566006 434898 566048 435134
rect 565728 434866 566048 434898
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 565728 399454 566048 399486
rect 565728 399218 565770 399454
rect 566006 399218 566048 399454
rect 565728 399134 566048 399218
rect 565728 398898 565770 399134
rect 566006 398898 566048 399134
rect 565728 398866 566048 398898
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 565728 363454 566048 363486
rect 565728 363218 565770 363454
rect 566006 363218 566048 363454
rect 565728 363134 566048 363218
rect 565728 362898 565770 363134
rect 566006 362898 566048 363134
rect 565728 362866 566048 362898
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 565728 327454 566048 327486
rect 565728 327218 565770 327454
rect 566006 327218 566048 327454
rect 565728 327134 566048 327218
rect 565728 326898 565770 327134
rect 566006 326898 566048 327134
rect 565728 326866 566048 326898
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 565728 291454 566048 291486
rect 565728 291218 565770 291454
rect 566006 291218 566048 291454
rect 565728 291134 566048 291218
rect 565728 290898 565770 291134
rect 566006 290898 566048 291134
rect 565728 290866 566048 290898
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 565728 255454 566048 255486
rect 565728 255218 565770 255454
rect 566006 255218 566048 255454
rect 565728 255134 566048 255218
rect 565728 254898 565770 255134
rect 566006 254898 566048 255134
rect 565728 254866 566048 254898
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 565728 219454 566048 219486
rect 565728 219218 565770 219454
rect 566006 219218 566048 219454
rect 565728 219134 566048 219218
rect 565728 218898 565770 219134
rect 566006 218898 566048 219134
rect 565728 218866 566048 218898
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 565728 183454 566048 183486
rect 565728 183218 565770 183454
rect 566006 183218 566048 183454
rect 565728 183134 566048 183218
rect 565728 182898 565770 183134
rect 566006 182898 566048 183134
rect 565728 182866 566048 182898
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 565728 147454 566048 147486
rect 565728 147218 565770 147454
rect 566006 147218 566048 147454
rect 565728 147134 566048 147218
rect 565728 146898 565770 147134
rect 566006 146898 566048 147134
rect 565728 146866 566048 146898
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 565728 111454 566048 111486
rect 565728 111218 565770 111454
rect 566006 111218 566048 111454
rect 565728 111134 566048 111218
rect 565728 110898 565770 111134
rect 566006 110898 566048 111134
rect 565728 110866 566048 110898
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 565728 75454 566048 75486
rect 565728 75218 565770 75454
rect 566006 75218 566048 75454
rect 565728 75134 566048 75218
rect 565728 74898 565770 75134
rect 566006 74898 566048 75134
rect 565728 74866 566048 74898
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 552954 50614 553574 66000
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 550771 4860 550837 4861
rect 550771 4796 550772 4860
rect 550836 4796 550837 4860
rect 550771 4795 550837 4796
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 57454 560414 66000
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 61174 564134 66000
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 64894 567854 66000
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 32614 571574 66000
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 74250 543218 74486 543454
rect 74250 542898 74486 543134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 74250 507218 74486 507454
rect 74250 506898 74486 507134
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 74250 471218 74486 471454
rect 74250 470898 74486 471134
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 74250 435218 74486 435454
rect 74250 434898 74486 435134
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 74250 399218 74486 399454
rect 74250 398898 74486 399134
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 74250 327218 74486 327454
rect 74250 326898 74486 327134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 74250 291218 74486 291454
rect 74250 290898 74486 291134
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 74250 219218 74486 219454
rect 74250 218898 74486 219134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 74250 183218 74486 183454
rect 74250 182898 74486 183134
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 74250 147218 74486 147454
rect 74250 146898 74486 147134
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 74250 111218 74486 111454
rect 74250 110898 74486 111134
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 74250 75218 74486 75454
rect 74250 74898 74486 75134
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 89610 561218 89846 561454
rect 89610 560898 89846 561134
rect 89610 525218 89846 525454
rect 89610 524898 89846 525134
rect 89610 489218 89846 489454
rect 89610 488898 89846 489134
rect 89610 453218 89846 453454
rect 89610 452898 89846 453134
rect 89610 417218 89846 417454
rect 89610 416898 89846 417134
rect 89610 381218 89846 381454
rect 89610 380898 89846 381134
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 89610 309218 89846 309454
rect 89610 308898 89846 309134
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 89610 237218 89846 237454
rect 89610 236898 89846 237134
rect 89610 201218 89846 201454
rect 89610 200898 89846 201134
rect 89610 165218 89846 165454
rect 89610 164898 89846 165134
rect 89610 129218 89846 129454
rect 89610 128898 89846 129134
rect 89610 93218 89846 93454
rect 89610 92898 89846 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 104970 543218 105206 543454
rect 104970 542898 105206 543134
rect 104970 507218 105206 507454
rect 104970 506898 105206 507134
rect 104970 471218 105206 471454
rect 104970 470898 105206 471134
rect 104970 435218 105206 435454
rect 104970 434898 105206 435134
rect 104970 399218 105206 399454
rect 104970 398898 105206 399134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 104970 327218 105206 327454
rect 104970 326898 105206 327134
rect 104970 291218 105206 291454
rect 104970 290898 105206 291134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 104970 219218 105206 219454
rect 104970 218898 105206 219134
rect 104970 183218 105206 183454
rect 104970 182898 105206 183134
rect 104970 147218 105206 147454
rect 104970 146898 105206 147134
rect 104970 111218 105206 111454
rect 104970 110898 105206 111134
rect 104970 75218 105206 75454
rect 104970 74898 105206 75134
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 120330 561218 120566 561454
rect 120330 560898 120566 561134
rect 120330 525218 120566 525454
rect 120330 524898 120566 525134
rect 120330 489218 120566 489454
rect 120330 488898 120566 489134
rect 120330 453218 120566 453454
rect 120330 452898 120566 453134
rect 120330 417218 120566 417454
rect 120330 416898 120566 417134
rect 120330 381218 120566 381454
rect 120330 380898 120566 381134
rect 120330 345218 120566 345454
rect 120330 344898 120566 345134
rect 120330 309218 120566 309454
rect 120330 308898 120566 309134
rect 120330 273218 120566 273454
rect 120330 272898 120566 273134
rect 120330 237218 120566 237454
rect 120330 236898 120566 237134
rect 120330 201218 120566 201454
rect 120330 200898 120566 201134
rect 120330 165218 120566 165454
rect 120330 164898 120566 165134
rect 120330 129218 120566 129454
rect 120330 128898 120566 129134
rect 120330 93218 120566 93454
rect 120330 92898 120566 93134
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 135690 543218 135926 543454
rect 135690 542898 135926 543134
rect 135690 507218 135926 507454
rect 135690 506898 135926 507134
rect 135690 471218 135926 471454
rect 135690 470898 135926 471134
rect 135690 435218 135926 435454
rect 135690 434898 135926 435134
rect 135690 399218 135926 399454
rect 135690 398898 135926 399134
rect 135690 363218 135926 363454
rect 135690 362898 135926 363134
rect 135690 327218 135926 327454
rect 135690 326898 135926 327134
rect 135690 291218 135926 291454
rect 135690 290898 135926 291134
rect 135690 255218 135926 255454
rect 135690 254898 135926 255134
rect 135690 219218 135926 219454
rect 135690 218898 135926 219134
rect 135690 183218 135926 183454
rect 135690 182898 135926 183134
rect 135690 147218 135926 147454
rect 135690 146898 135926 147134
rect 135690 111218 135926 111454
rect 135690 110898 135926 111134
rect 135690 75218 135926 75454
rect 135690 74898 135926 75134
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 151050 561218 151286 561454
rect 151050 560898 151286 561134
rect 151050 525218 151286 525454
rect 151050 524898 151286 525134
rect 151050 489218 151286 489454
rect 151050 488898 151286 489134
rect 151050 453218 151286 453454
rect 151050 452898 151286 453134
rect 151050 417218 151286 417454
rect 151050 416898 151286 417134
rect 151050 381218 151286 381454
rect 151050 380898 151286 381134
rect 151050 345218 151286 345454
rect 151050 344898 151286 345134
rect 151050 309218 151286 309454
rect 151050 308898 151286 309134
rect 151050 273218 151286 273454
rect 151050 272898 151286 273134
rect 151050 237218 151286 237454
rect 151050 236898 151286 237134
rect 151050 201218 151286 201454
rect 151050 200898 151286 201134
rect 151050 165218 151286 165454
rect 151050 164898 151286 165134
rect 151050 129218 151286 129454
rect 151050 128898 151286 129134
rect 151050 93218 151286 93454
rect 151050 92898 151286 93134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 166410 543218 166646 543454
rect 166410 542898 166646 543134
rect 166410 507218 166646 507454
rect 166410 506898 166646 507134
rect 166410 471218 166646 471454
rect 166410 470898 166646 471134
rect 166410 435218 166646 435454
rect 166410 434898 166646 435134
rect 166410 399218 166646 399454
rect 166410 398898 166646 399134
rect 166410 363218 166646 363454
rect 166410 362898 166646 363134
rect 166410 327218 166646 327454
rect 166410 326898 166646 327134
rect 166410 291218 166646 291454
rect 166410 290898 166646 291134
rect 166410 255218 166646 255454
rect 166410 254898 166646 255134
rect 166410 219218 166646 219454
rect 166410 218898 166646 219134
rect 166410 183218 166646 183454
rect 166410 182898 166646 183134
rect 166410 147218 166646 147454
rect 166410 146898 166646 147134
rect 166410 111218 166646 111454
rect 166410 110898 166646 111134
rect 166410 75218 166646 75454
rect 166410 74898 166646 75134
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 181770 561218 182006 561454
rect 181770 560898 182006 561134
rect 197130 543218 197366 543454
rect 197130 542898 197366 543134
rect 181770 525218 182006 525454
rect 181770 524898 182006 525134
rect 197130 507218 197366 507454
rect 197130 506898 197366 507134
rect 181770 489218 182006 489454
rect 181770 488898 182006 489134
rect 197130 471218 197366 471454
rect 197130 470898 197366 471134
rect 181770 453218 182006 453454
rect 181770 452898 182006 453134
rect 197130 435218 197366 435454
rect 197130 434898 197366 435134
rect 181770 417218 182006 417454
rect 181770 416898 182006 417134
rect 197130 399218 197366 399454
rect 197130 398898 197366 399134
rect 181770 381218 182006 381454
rect 181770 380898 182006 381134
rect 197130 363218 197366 363454
rect 197130 362898 197366 363134
rect 181770 345218 182006 345454
rect 181770 344898 182006 345134
rect 197130 327218 197366 327454
rect 197130 326898 197366 327134
rect 181770 309218 182006 309454
rect 181770 308898 182006 309134
rect 197130 291218 197366 291454
rect 197130 290898 197366 291134
rect 181770 273218 182006 273454
rect 181770 272898 182006 273134
rect 197130 255218 197366 255454
rect 197130 254898 197366 255134
rect 181770 237218 182006 237454
rect 181770 236898 182006 237134
rect 197130 219218 197366 219454
rect 197130 218898 197366 219134
rect 181770 201218 182006 201454
rect 181770 200898 182006 201134
rect 197130 183218 197366 183454
rect 197130 182898 197366 183134
rect 181770 165218 182006 165454
rect 181770 164898 182006 165134
rect 197130 147218 197366 147454
rect 197130 146898 197366 147134
rect 181770 129218 182006 129454
rect 181770 128898 182006 129134
rect 197130 111218 197366 111454
rect 197130 110898 197366 111134
rect 181770 93218 182006 93454
rect 181770 92898 182006 93134
rect 197130 75218 197366 75454
rect 197130 74898 197366 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 212490 561218 212726 561454
rect 212490 560898 212726 561134
rect 212490 525218 212726 525454
rect 212490 524898 212726 525134
rect 212490 489218 212726 489454
rect 212490 488898 212726 489134
rect 212490 453218 212726 453454
rect 212490 452898 212726 453134
rect 212490 417218 212726 417454
rect 212490 416898 212726 417134
rect 212490 381218 212726 381454
rect 212490 380898 212726 381134
rect 212490 345218 212726 345454
rect 212490 344898 212726 345134
rect 212490 309218 212726 309454
rect 212490 308898 212726 309134
rect 212490 273218 212726 273454
rect 212490 272898 212726 273134
rect 212490 237218 212726 237454
rect 212490 236898 212726 237134
rect 212490 201218 212726 201454
rect 212490 200898 212726 201134
rect 212490 165218 212726 165454
rect 212490 164898 212726 165134
rect 212490 129218 212726 129454
rect 212490 128898 212726 129134
rect 212490 93218 212726 93454
rect 212490 92898 212726 93134
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 227850 543218 228086 543454
rect 227850 542898 228086 543134
rect 227850 507218 228086 507454
rect 227850 506898 228086 507134
rect 227850 471218 228086 471454
rect 227850 470898 228086 471134
rect 227850 435218 228086 435454
rect 227850 434898 228086 435134
rect 227850 399218 228086 399454
rect 227850 398898 228086 399134
rect 227850 363218 228086 363454
rect 227850 362898 228086 363134
rect 227850 327218 228086 327454
rect 227850 326898 228086 327134
rect 227850 291218 228086 291454
rect 227850 290898 228086 291134
rect 227850 255218 228086 255454
rect 227850 254898 228086 255134
rect 227850 219218 228086 219454
rect 227850 218898 228086 219134
rect 227850 183218 228086 183454
rect 227850 182898 228086 183134
rect 227850 147218 228086 147454
rect 227850 146898 228086 147134
rect 227850 111218 228086 111454
rect 227850 110898 228086 111134
rect 227850 75218 228086 75454
rect 227850 74898 228086 75134
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 243210 561218 243446 561454
rect 243210 560898 243446 561134
rect 243210 525218 243446 525454
rect 243210 524898 243446 525134
rect 243210 489218 243446 489454
rect 243210 488898 243446 489134
rect 243210 453218 243446 453454
rect 243210 452898 243446 453134
rect 243210 417218 243446 417454
rect 243210 416898 243446 417134
rect 243210 381218 243446 381454
rect 243210 380898 243446 381134
rect 243210 345218 243446 345454
rect 243210 344898 243446 345134
rect 243210 309218 243446 309454
rect 243210 308898 243446 309134
rect 243210 273218 243446 273454
rect 243210 272898 243446 273134
rect 243210 237218 243446 237454
rect 243210 236898 243446 237134
rect 243210 201218 243446 201454
rect 243210 200898 243446 201134
rect 243210 165218 243446 165454
rect 243210 164898 243446 165134
rect 243210 129218 243446 129454
rect 243210 128898 243446 129134
rect 243210 93218 243446 93454
rect 243210 92898 243446 93134
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 258570 543218 258806 543454
rect 258570 542898 258806 543134
rect 258570 507218 258806 507454
rect 258570 506898 258806 507134
rect 258570 471218 258806 471454
rect 258570 470898 258806 471134
rect 258570 435218 258806 435454
rect 258570 434898 258806 435134
rect 258570 399218 258806 399454
rect 258570 398898 258806 399134
rect 258570 363218 258806 363454
rect 258570 362898 258806 363134
rect 258570 327218 258806 327454
rect 258570 326898 258806 327134
rect 258570 291218 258806 291454
rect 258570 290898 258806 291134
rect 258570 255218 258806 255454
rect 258570 254898 258806 255134
rect 258570 219218 258806 219454
rect 258570 218898 258806 219134
rect 258570 183218 258806 183454
rect 258570 182898 258806 183134
rect 258570 147218 258806 147454
rect 258570 146898 258806 147134
rect 258570 111218 258806 111454
rect 258570 110898 258806 111134
rect 258570 75218 258806 75454
rect 258570 74898 258806 75134
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 273930 561218 274166 561454
rect 273930 560898 274166 561134
rect 273930 525218 274166 525454
rect 273930 524898 274166 525134
rect 273930 489218 274166 489454
rect 273930 488898 274166 489134
rect 273930 453218 274166 453454
rect 273930 452898 274166 453134
rect 273930 417218 274166 417454
rect 273930 416898 274166 417134
rect 273930 381218 274166 381454
rect 273930 380898 274166 381134
rect 273930 345218 274166 345454
rect 273930 344898 274166 345134
rect 273930 309218 274166 309454
rect 273930 308898 274166 309134
rect 273930 273218 274166 273454
rect 273930 272898 274166 273134
rect 273930 237218 274166 237454
rect 273930 236898 274166 237134
rect 273930 201218 274166 201454
rect 273930 200898 274166 201134
rect 273930 165218 274166 165454
rect 273930 164898 274166 165134
rect 273930 129218 274166 129454
rect 273930 128898 274166 129134
rect 273930 93218 274166 93454
rect 273930 92898 274166 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 304650 561218 304886 561454
rect 304650 560898 304886 561134
rect 335370 561218 335606 561454
rect 335370 560898 335606 561134
rect 289290 543218 289526 543454
rect 289290 542898 289526 543134
rect 320010 543218 320246 543454
rect 320010 542898 320246 543134
rect 304650 525218 304886 525454
rect 304650 524898 304886 525134
rect 335370 525218 335606 525454
rect 335370 524898 335606 525134
rect 289290 507218 289526 507454
rect 289290 506898 289526 507134
rect 320010 507218 320246 507454
rect 320010 506898 320246 507134
rect 304650 489218 304886 489454
rect 304650 488898 304886 489134
rect 335370 489218 335606 489454
rect 335370 488898 335606 489134
rect 289290 471218 289526 471454
rect 289290 470898 289526 471134
rect 320010 471218 320246 471454
rect 320010 470898 320246 471134
rect 304650 453218 304886 453454
rect 304650 452898 304886 453134
rect 335370 453218 335606 453454
rect 335370 452898 335606 453134
rect 289290 435218 289526 435454
rect 289290 434898 289526 435134
rect 320010 435218 320246 435454
rect 320010 434898 320246 435134
rect 304650 417218 304886 417454
rect 304650 416898 304886 417134
rect 335370 417218 335606 417454
rect 335370 416898 335606 417134
rect 289290 399218 289526 399454
rect 289290 398898 289526 399134
rect 320010 399218 320246 399454
rect 320010 398898 320246 399134
rect 304650 381218 304886 381454
rect 304650 380898 304886 381134
rect 335370 381218 335606 381454
rect 335370 380898 335606 381134
rect 289290 363218 289526 363454
rect 289290 362898 289526 363134
rect 320010 363218 320246 363454
rect 320010 362898 320246 363134
rect 304650 345218 304886 345454
rect 304650 344898 304886 345134
rect 335370 345218 335606 345454
rect 335370 344898 335606 345134
rect 289290 327218 289526 327454
rect 289290 326898 289526 327134
rect 320010 327218 320246 327454
rect 320010 326898 320246 327134
rect 304650 309218 304886 309454
rect 304650 308898 304886 309134
rect 335370 309218 335606 309454
rect 335370 308898 335606 309134
rect 289290 291218 289526 291454
rect 289290 290898 289526 291134
rect 320010 291218 320246 291454
rect 320010 290898 320246 291134
rect 304650 273218 304886 273454
rect 304650 272898 304886 273134
rect 335370 273218 335606 273454
rect 335370 272898 335606 273134
rect 289290 255218 289526 255454
rect 289290 254898 289526 255134
rect 320010 255218 320246 255454
rect 320010 254898 320246 255134
rect 304650 237218 304886 237454
rect 304650 236898 304886 237134
rect 335370 237218 335606 237454
rect 335370 236898 335606 237134
rect 289290 219218 289526 219454
rect 289290 218898 289526 219134
rect 320010 219218 320246 219454
rect 320010 218898 320246 219134
rect 304650 201218 304886 201454
rect 304650 200898 304886 201134
rect 335370 201218 335606 201454
rect 335370 200898 335606 201134
rect 289290 183218 289526 183454
rect 289290 182898 289526 183134
rect 320010 183218 320246 183454
rect 320010 182898 320246 183134
rect 304650 165218 304886 165454
rect 304650 164898 304886 165134
rect 335370 165218 335606 165454
rect 335370 164898 335606 165134
rect 289290 147218 289526 147454
rect 289290 146898 289526 147134
rect 320010 147218 320246 147454
rect 320010 146898 320246 147134
rect 304650 129218 304886 129454
rect 304650 128898 304886 129134
rect 335370 129218 335606 129454
rect 335370 128898 335606 129134
rect 289290 111218 289526 111454
rect 289290 110898 289526 111134
rect 320010 111218 320246 111454
rect 320010 110898 320246 111134
rect 304650 93218 304886 93454
rect 304650 92898 304886 93134
rect 335370 93218 335606 93454
rect 335370 92898 335606 93134
rect 289290 75218 289526 75454
rect 289290 74898 289526 75134
rect 320010 75218 320246 75454
rect 320010 74898 320246 75134
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 366090 561218 366326 561454
rect 366090 560898 366326 561134
rect 350730 543218 350966 543454
rect 350730 542898 350966 543134
rect 381450 543218 381686 543454
rect 381450 542898 381686 543134
rect 366090 525218 366326 525454
rect 366090 524898 366326 525134
rect 350730 507218 350966 507454
rect 350730 506898 350966 507134
rect 381450 507218 381686 507454
rect 381450 506898 381686 507134
rect 366090 489218 366326 489454
rect 366090 488898 366326 489134
rect 350730 471218 350966 471454
rect 350730 470898 350966 471134
rect 381450 471218 381686 471454
rect 381450 470898 381686 471134
rect 366090 453218 366326 453454
rect 366090 452898 366326 453134
rect 350730 435218 350966 435454
rect 350730 434898 350966 435134
rect 381450 435218 381686 435454
rect 381450 434898 381686 435134
rect 366090 417218 366326 417454
rect 366090 416898 366326 417134
rect 350730 399218 350966 399454
rect 350730 398898 350966 399134
rect 381450 399218 381686 399454
rect 381450 398898 381686 399134
rect 366090 381218 366326 381454
rect 366090 380898 366326 381134
rect 350730 363218 350966 363454
rect 350730 362898 350966 363134
rect 381450 363218 381686 363454
rect 381450 362898 381686 363134
rect 366090 345218 366326 345454
rect 366090 344898 366326 345134
rect 350730 327218 350966 327454
rect 350730 326898 350966 327134
rect 381450 327218 381686 327454
rect 381450 326898 381686 327134
rect 366090 309218 366326 309454
rect 366090 308898 366326 309134
rect 350730 291218 350966 291454
rect 350730 290898 350966 291134
rect 381450 291218 381686 291454
rect 381450 290898 381686 291134
rect 366090 273218 366326 273454
rect 366090 272898 366326 273134
rect 350730 255218 350966 255454
rect 350730 254898 350966 255134
rect 381450 255218 381686 255454
rect 381450 254898 381686 255134
rect 366090 237218 366326 237454
rect 366090 236898 366326 237134
rect 350730 219218 350966 219454
rect 350730 218898 350966 219134
rect 381450 219218 381686 219454
rect 381450 218898 381686 219134
rect 366090 201218 366326 201454
rect 366090 200898 366326 201134
rect 350730 183218 350966 183454
rect 350730 182898 350966 183134
rect 381450 183218 381686 183454
rect 381450 182898 381686 183134
rect 366090 165218 366326 165454
rect 366090 164898 366326 165134
rect 350730 147218 350966 147454
rect 350730 146898 350966 147134
rect 381450 147218 381686 147454
rect 381450 146898 381686 147134
rect 366090 129218 366326 129454
rect 366090 128898 366326 129134
rect 350730 111218 350966 111454
rect 350730 110898 350966 111134
rect 381450 111218 381686 111454
rect 381450 110898 381686 111134
rect 366090 93218 366326 93454
rect 366090 92898 366326 93134
rect 350730 75218 350966 75454
rect 350730 74898 350966 75134
rect 381450 75218 381686 75454
rect 381450 74898 381686 75134
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 396810 561218 397046 561454
rect 396810 560898 397046 561134
rect 396810 525218 397046 525454
rect 396810 524898 397046 525134
rect 396810 489218 397046 489454
rect 396810 488898 397046 489134
rect 396810 453218 397046 453454
rect 396810 452898 397046 453134
rect 396810 417218 397046 417454
rect 396810 416898 397046 417134
rect 396810 381218 397046 381454
rect 396810 380898 397046 381134
rect 396810 345218 397046 345454
rect 396810 344898 397046 345134
rect 396810 309218 397046 309454
rect 396810 308898 397046 309134
rect 396810 273218 397046 273454
rect 396810 272898 397046 273134
rect 396810 237218 397046 237454
rect 396810 236898 397046 237134
rect 396810 201218 397046 201454
rect 396810 200898 397046 201134
rect 396810 165218 397046 165454
rect 396810 164898 397046 165134
rect 396810 129218 397046 129454
rect 396810 128898 397046 129134
rect 396810 93218 397046 93454
rect 396810 92898 397046 93134
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 427530 561218 427766 561454
rect 427530 560898 427766 561134
rect 412170 543218 412406 543454
rect 412170 542898 412406 543134
rect 427530 525218 427766 525454
rect 427530 524898 427766 525134
rect 412170 507218 412406 507454
rect 412170 506898 412406 507134
rect 427530 489218 427766 489454
rect 427530 488898 427766 489134
rect 412170 471218 412406 471454
rect 412170 470898 412406 471134
rect 427530 453218 427766 453454
rect 427530 452898 427766 453134
rect 412170 435218 412406 435454
rect 412170 434898 412406 435134
rect 427530 417218 427766 417454
rect 427530 416898 427766 417134
rect 412170 399218 412406 399454
rect 412170 398898 412406 399134
rect 427530 381218 427766 381454
rect 427530 380898 427766 381134
rect 412170 363218 412406 363454
rect 412170 362898 412406 363134
rect 427530 345218 427766 345454
rect 427530 344898 427766 345134
rect 412170 327218 412406 327454
rect 412170 326898 412406 327134
rect 427530 309218 427766 309454
rect 427530 308898 427766 309134
rect 412170 291218 412406 291454
rect 412170 290898 412406 291134
rect 427530 273218 427766 273454
rect 427530 272898 427766 273134
rect 412170 255218 412406 255454
rect 412170 254898 412406 255134
rect 427530 237218 427766 237454
rect 427530 236898 427766 237134
rect 412170 219218 412406 219454
rect 412170 218898 412406 219134
rect 427530 201218 427766 201454
rect 427530 200898 427766 201134
rect 412170 183218 412406 183454
rect 412170 182898 412406 183134
rect 427530 165218 427766 165454
rect 427530 164898 427766 165134
rect 412170 147218 412406 147454
rect 412170 146898 412406 147134
rect 427530 129218 427766 129454
rect 427530 128898 427766 129134
rect 412170 111218 412406 111454
rect 412170 110898 412406 111134
rect 427530 93218 427766 93454
rect 427530 92898 427766 93134
rect 412170 75218 412406 75454
rect 412170 74898 412406 75134
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 458250 561218 458486 561454
rect 458250 560898 458486 561134
rect 442890 543218 443126 543454
rect 442890 542898 443126 543134
rect 458250 525218 458486 525454
rect 458250 524898 458486 525134
rect 442890 507218 443126 507454
rect 442890 506898 443126 507134
rect 458250 489218 458486 489454
rect 458250 488898 458486 489134
rect 442890 471218 443126 471454
rect 442890 470898 443126 471134
rect 458250 453218 458486 453454
rect 458250 452898 458486 453134
rect 442890 435218 443126 435454
rect 442890 434898 443126 435134
rect 458250 417218 458486 417454
rect 458250 416898 458486 417134
rect 442890 399218 443126 399454
rect 442890 398898 443126 399134
rect 458250 381218 458486 381454
rect 458250 380898 458486 381134
rect 442890 363218 443126 363454
rect 442890 362898 443126 363134
rect 458250 345218 458486 345454
rect 458250 344898 458486 345134
rect 442890 327218 443126 327454
rect 442890 326898 443126 327134
rect 458250 309218 458486 309454
rect 458250 308898 458486 309134
rect 442890 291218 443126 291454
rect 442890 290898 443126 291134
rect 458250 273218 458486 273454
rect 458250 272898 458486 273134
rect 442890 255218 443126 255454
rect 442890 254898 443126 255134
rect 458250 237218 458486 237454
rect 458250 236898 458486 237134
rect 442890 219218 443126 219454
rect 442890 218898 443126 219134
rect 458250 201218 458486 201454
rect 458250 200898 458486 201134
rect 442890 183218 443126 183454
rect 442890 182898 443126 183134
rect 458250 165218 458486 165454
rect 458250 164898 458486 165134
rect 442890 147218 443126 147454
rect 442890 146898 443126 147134
rect 458250 129218 458486 129454
rect 458250 128898 458486 129134
rect 442890 111218 443126 111454
rect 442890 110898 443126 111134
rect 458250 93218 458486 93454
rect 458250 92898 458486 93134
rect 442890 75218 443126 75454
rect 442890 74898 443126 75134
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 473610 543218 473846 543454
rect 473610 542898 473846 543134
rect 473610 507218 473846 507454
rect 473610 506898 473846 507134
rect 473610 471218 473846 471454
rect 473610 470898 473846 471134
rect 473610 435218 473846 435454
rect 473610 434898 473846 435134
rect 473610 399218 473846 399454
rect 473610 398898 473846 399134
rect 473610 363218 473846 363454
rect 473610 362898 473846 363134
rect 473610 327218 473846 327454
rect 473610 326898 473846 327134
rect 473610 291218 473846 291454
rect 473610 290898 473846 291134
rect 473610 255218 473846 255454
rect 473610 254898 473846 255134
rect 473610 219218 473846 219454
rect 473610 218898 473846 219134
rect 473610 183218 473846 183454
rect 473610 182898 473846 183134
rect 473610 147218 473846 147454
rect 473610 146898 473846 147134
rect 473610 111218 473846 111454
rect 473610 110898 473846 111134
rect 473610 75218 473846 75454
rect 473610 74898 473846 75134
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 488970 561218 489206 561454
rect 488970 560898 489206 561134
rect 519690 561218 519926 561454
rect 519690 560898 519926 561134
rect 504330 543218 504566 543454
rect 504330 542898 504566 543134
rect 535050 543218 535286 543454
rect 535050 542898 535286 543134
rect 488970 525218 489206 525454
rect 488970 524898 489206 525134
rect 519690 525218 519926 525454
rect 519690 524898 519926 525134
rect 504330 507218 504566 507454
rect 504330 506898 504566 507134
rect 535050 507218 535286 507454
rect 535050 506898 535286 507134
rect 488970 489218 489206 489454
rect 488970 488898 489206 489134
rect 519690 489218 519926 489454
rect 519690 488898 519926 489134
rect 504330 471218 504566 471454
rect 504330 470898 504566 471134
rect 535050 471218 535286 471454
rect 535050 470898 535286 471134
rect 488970 453218 489206 453454
rect 488970 452898 489206 453134
rect 519690 453218 519926 453454
rect 519690 452898 519926 453134
rect 504330 435218 504566 435454
rect 504330 434898 504566 435134
rect 535050 435218 535286 435454
rect 535050 434898 535286 435134
rect 488970 417218 489206 417454
rect 488970 416898 489206 417134
rect 519690 417218 519926 417454
rect 519690 416898 519926 417134
rect 504330 399218 504566 399454
rect 504330 398898 504566 399134
rect 535050 399218 535286 399454
rect 535050 398898 535286 399134
rect 488970 381218 489206 381454
rect 488970 380898 489206 381134
rect 519690 381218 519926 381454
rect 519690 380898 519926 381134
rect 504330 363218 504566 363454
rect 504330 362898 504566 363134
rect 535050 363218 535286 363454
rect 535050 362898 535286 363134
rect 488970 345218 489206 345454
rect 488970 344898 489206 345134
rect 519690 345218 519926 345454
rect 519690 344898 519926 345134
rect 504330 327218 504566 327454
rect 504330 326898 504566 327134
rect 535050 327218 535286 327454
rect 535050 326898 535286 327134
rect 488970 309218 489206 309454
rect 488970 308898 489206 309134
rect 519690 309218 519926 309454
rect 519690 308898 519926 309134
rect 504330 291218 504566 291454
rect 504330 290898 504566 291134
rect 535050 291218 535286 291454
rect 535050 290898 535286 291134
rect 488970 273218 489206 273454
rect 488970 272898 489206 273134
rect 519690 273218 519926 273454
rect 519690 272898 519926 273134
rect 504330 255218 504566 255454
rect 504330 254898 504566 255134
rect 535050 255218 535286 255454
rect 535050 254898 535286 255134
rect 488970 237218 489206 237454
rect 488970 236898 489206 237134
rect 519690 237218 519926 237454
rect 519690 236898 519926 237134
rect 504330 219218 504566 219454
rect 504330 218898 504566 219134
rect 535050 219218 535286 219454
rect 535050 218898 535286 219134
rect 488970 201218 489206 201454
rect 488970 200898 489206 201134
rect 519690 201218 519926 201454
rect 519690 200898 519926 201134
rect 504330 183218 504566 183454
rect 504330 182898 504566 183134
rect 535050 183218 535286 183454
rect 535050 182898 535286 183134
rect 488970 165218 489206 165454
rect 488970 164898 489206 165134
rect 519690 165218 519926 165454
rect 519690 164898 519926 165134
rect 504330 147218 504566 147454
rect 504330 146898 504566 147134
rect 535050 147218 535286 147454
rect 535050 146898 535286 147134
rect 488970 129218 489206 129454
rect 488970 128898 489206 129134
rect 519690 129218 519926 129454
rect 519690 128898 519926 129134
rect 504330 111218 504566 111454
rect 504330 110898 504566 111134
rect 535050 111218 535286 111454
rect 535050 110898 535286 111134
rect 488970 93218 489206 93454
rect 488970 92898 489206 93134
rect 519690 93218 519926 93454
rect 519690 92898 519926 93134
rect 504330 75218 504566 75454
rect 504330 74898 504566 75134
rect 535050 75218 535286 75454
rect 535050 74898 535286 75134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 550410 561218 550646 561454
rect 550410 560898 550646 561134
rect 550410 525218 550646 525454
rect 550410 524898 550646 525134
rect 550410 489218 550646 489454
rect 550410 488898 550646 489134
rect 550410 453218 550646 453454
rect 550410 452898 550646 453134
rect 550410 417218 550646 417454
rect 550410 416898 550646 417134
rect 550410 381218 550646 381454
rect 550410 380898 550646 381134
rect 550410 345218 550646 345454
rect 550410 344898 550646 345134
rect 550410 309218 550646 309454
rect 550410 308898 550646 309134
rect 550410 273218 550646 273454
rect 550410 272898 550646 273134
rect 550410 237218 550646 237454
rect 550410 236898 550646 237134
rect 550410 201218 550646 201454
rect 550410 200898 550646 201134
rect 550410 165218 550646 165454
rect 550410 164898 550646 165134
rect 550410 129218 550646 129454
rect 550410 128898 550646 129134
rect 550410 93218 550646 93454
rect 550410 92898 550646 93134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 565770 543218 566006 543454
rect 565770 542898 566006 543134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 565770 507218 566006 507454
rect 565770 506898 566006 507134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 565770 471218 566006 471454
rect 565770 470898 566006 471134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 565770 435218 566006 435454
rect 565770 434898 566006 435134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 565770 399218 566006 399454
rect 565770 398898 566006 399134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 565770 363218 566006 363454
rect 565770 362898 566006 363134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 565770 327218 566006 327454
rect 565770 326898 566006 327134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 565770 291218 566006 291454
rect 565770 290898 566006 291134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 565770 255218 566006 255454
rect 565770 254898 566006 255134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 565770 219218 566006 219454
rect 565770 218898 566006 219134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 565770 183218 566006 183454
rect 565770 182898 566006 183134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 565770 147218 566006 147454
rect 565770 146898 566006 147134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 565770 111218 566006 111454
rect 565770 110898 566006 111134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 565770 75218 566006 75454
rect 565770 74898 566006 75134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 89610 561454
rect 89846 561218 120330 561454
rect 120566 561218 151050 561454
rect 151286 561218 181770 561454
rect 182006 561218 212490 561454
rect 212726 561218 243210 561454
rect 243446 561218 273930 561454
rect 274166 561218 304650 561454
rect 304886 561218 335370 561454
rect 335606 561218 366090 561454
rect 366326 561218 396810 561454
rect 397046 561218 427530 561454
rect 427766 561218 458250 561454
rect 458486 561218 488970 561454
rect 489206 561218 519690 561454
rect 519926 561218 550410 561454
rect 550646 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 89610 561134
rect 89846 560898 120330 561134
rect 120566 560898 151050 561134
rect 151286 560898 181770 561134
rect 182006 560898 212490 561134
rect 212726 560898 243210 561134
rect 243446 560898 273930 561134
rect 274166 560898 304650 561134
rect 304886 560898 335370 561134
rect 335606 560898 366090 561134
rect 366326 560898 396810 561134
rect 397046 560898 427530 561134
rect 427766 560898 458250 561134
rect 458486 560898 488970 561134
rect 489206 560898 519690 561134
rect 519926 560898 550410 561134
rect 550646 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 74250 543454
rect 74486 543218 104970 543454
rect 105206 543218 135690 543454
rect 135926 543218 166410 543454
rect 166646 543218 197130 543454
rect 197366 543218 227850 543454
rect 228086 543218 258570 543454
rect 258806 543218 289290 543454
rect 289526 543218 320010 543454
rect 320246 543218 350730 543454
rect 350966 543218 381450 543454
rect 381686 543218 412170 543454
rect 412406 543218 442890 543454
rect 443126 543218 473610 543454
rect 473846 543218 504330 543454
rect 504566 543218 535050 543454
rect 535286 543218 565770 543454
rect 566006 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 74250 543134
rect 74486 542898 104970 543134
rect 105206 542898 135690 543134
rect 135926 542898 166410 543134
rect 166646 542898 197130 543134
rect 197366 542898 227850 543134
rect 228086 542898 258570 543134
rect 258806 542898 289290 543134
rect 289526 542898 320010 543134
rect 320246 542898 350730 543134
rect 350966 542898 381450 543134
rect 381686 542898 412170 543134
rect 412406 542898 442890 543134
rect 443126 542898 473610 543134
rect 473846 542898 504330 543134
rect 504566 542898 535050 543134
rect 535286 542898 565770 543134
rect 566006 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 89610 525454
rect 89846 525218 120330 525454
rect 120566 525218 151050 525454
rect 151286 525218 181770 525454
rect 182006 525218 212490 525454
rect 212726 525218 243210 525454
rect 243446 525218 273930 525454
rect 274166 525218 304650 525454
rect 304886 525218 335370 525454
rect 335606 525218 366090 525454
rect 366326 525218 396810 525454
rect 397046 525218 427530 525454
rect 427766 525218 458250 525454
rect 458486 525218 488970 525454
rect 489206 525218 519690 525454
rect 519926 525218 550410 525454
rect 550646 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 89610 525134
rect 89846 524898 120330 525134
rect 120566 524898 151050 525134
rect 151286 524898 181770 525134
rect 182006 524898 212490 525134
rect 212726 524898 243210 525134
rect 243446 524898 273930 525134
rect 274166 524898 304650 525134
rect 304886 524898 335370 525134
rect 335606 524898 366090 525134
rect 366326 524898 396810 525134
rect 397046 524898 427530 525134
rect 427766 524898 458250 525134
rect 458486 524898 488970 525134
rect 489206 524898 519690 525134
rect 519926 524898 550410 525134
rect 550646 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 74250 507454
rect 74486 507218 104970 507454
rect 105206 507218 135690 507454
rect 135926 507218 166410 507454
rect 166646 507218 197130 507454
rect 197366 507218 227850 507454
rect 228086 507218 258570 507454
rect 258806 507218 289290 507454
rect 289526 507218 320010 507454
rect 320246 507218 350730 507454
rect 350966 507218 381450 507454
rect 381686 507218 412170 507454
rect 412406 507218 442890 507454
rect 443126 507218 473610 507454
rect 473846 507218 504330 507454
rect 504566 507218 535050 507454
rect 535286 507218 565770 507454
rect 566006 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 74250 507134
rect 74486 506898 104970 507134
rect 105206 506898 135690 507134
rect 135926 506898 166410 507134
rect 166646 506898 197130 507134
rect 197366 506898 227850 507134
rect 228086 506898 258570 507134
rect 258806 506898 289290 507134
rect 289526 506898 320010 507134
rect 320246 506898 350730 507134
rect 350966 506898 381450 507134
rect 381686 506898 412170 507134
rect 412406 506898 442890 507134
rect 443126 506898 473610 507134
rect 473846 506898 504330 507134
rect 504566 506898 535050 507134
rect 535286 506898 565770 507134
rect 566006 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 89610 489454
rect 89846 489218 120330 489454
rect 120566 489218 151050 489454
rect 151286 489218 181770 489454
rect 182006 489218 212490 489454
rect 212726 489218 243210 489454
rect 243446 489218 273930 489454
rect 274166 489218 304650 489454
rect 304886 489218 335370 489454
rect 335606 489218 366090 489454
rect 366326 489218 396810 489454
rect 397046 489218 427530 489454
rect 427766 489218 458250 489454
rect 458486 489218 488970 489454
rect 489206 489218 519690 489454
rect 519926 489218 550410 489454
rect 550646 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 89610 489134
rect 89846 488898 120330 489134
rect 120566 488898 151050 489134
rect 151286 488898 181770 489134
rect 182006 488898 212490 489134
rect 212726 488898 243210 489134
rect 243446 488898 273930 489134
rect 274166 488898 304650 489134
rect 304886 488898 335370 489134
rect 335606 488898 366090 489134
rect 366326 488898 396810 489134
rect 397046 488898 427530 489134
rect 427766 488898 458250 489134
rect 458486 488898 488970 489134
rect 489206 488898 519690 489134
rect 519926 488898 550410 489134
rect 550646 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 74250 471454
rect 74486 471218 104970 471454
rect 105206 471218 135690 471454
rect 135926 471218 166410 471454
rect 166646 471218 197130 471454
rect 197366 471218 227850 471454
rect 228086 471218 258570 471454
rect 258806 471218 289290 471454
rect 289526 471218 320010 471454
rect 320246 471218 350730 471454
rect 350966 471218 381450 471454
rect 381686 471218 412170 471454
rect 412406 471218 442890 471454
rect 443126 471218 473610 471454
rect 473846 471218 504330 471454
rect 504566 471218 535050 471454
rect 535286 471218 565770 471454
rect 566006 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 74250 471134
rect 74486 470898 104970 471134
rect 105206 470898 135690 471134
rect 135926 470898 166410 471134
rect 166646 470898 197130 471134
rect 197366 470898 227850 471134
rect 228086 470898 258570 471134
rect 258806 470898 289290 471134
rect 289526 470898 320010 471134
rect 320246 470898 350730 471134
rect 350966 470898 381450 471134
rect 381686 470898 412170 471134
rect 412406 470898 442890 471134
rect 443126 470898 473610 471134
rect 473846 470898 504330 471134
rect 504566 470898 535050 471134
rect 535286 470898 565770 471134
rect 566006 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 89610 453454
rect 89846 453218 120330 453454
rect 120566 453218 151050 453454
rect 151286 453218 181770 453454
rect 182006 453218 212490 453454
rect 212726 453218 243210 453454
rect 243446 453218 273930 453454
rect 274166 453218 304650 453454
rect 304886 453218 335370 453454
rect 335606 453218 366090 453454
rect 366326 453218 396810 453454
rect 397046 453218 427530 453454
rect 427766 453218 458250 453454
rect 458486 453218 488970 453454
rect 489206 453218 519690 453454
rect 519926 453218 550410 453454
rect 550646 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 89610 453134
rect 89846 452898 120330 453134
rect 120566 452898 151050 453134
rect 151286 452898 181770 453134
rect 182006 452898 212490 453134
rect 212726 452898 243210 453134
rect 243446 452898 273930 453134
rect 274166 452898 304650 453134
rect 304886 452898 335370 453134
rect 335606 452898 366090 453134
rect 366326 452898 396810 453134
rect 397046 452898 427530 453134
rect 427766 452898 458250 453134
rect 458486 452898 488970 453134
rect 489206 452898 519690 453134
rect 519926 452898 550410 453134
rect 550646 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 74250 435454
rect 74486 435218 104970 435454
rect 105206 435218 135690 435454
rect 135926 435218 166410 435454
rect 166646 435218 197130 435454
rect 197366 435218 227850 435454
rect 228086 435218 258570 435454
rect 258806 435218 289290 435454
rect 289526 435218 320010 435454
rect 320246 435218 350730 435454
rect 350966 435218 381450 435454
rect 381686 435218 412170 435454
rect 412406 435218 442890 435454
rect 443126 435218 473610 435454
rect 473846 435218 504330 435454
rect 504566 435218 535050 435454
rect 535286 435218 565770 435454
rect 566006 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 74250 435134
rect 74486 434898 104970 435134
rect 105206 434898 135690 435134
rect 135926 434898 166410 435134
rect 166646 434898 197130 435134
rect 197366 434898 227850 435134
rect 228086 434898 258570 435134
rect 258806 434898 289290 435134
rect 289526 434898 320010 435134
rect 320246 434898 350730 435134
rect 350966 434898 381450 435134
rect 381686 434898 412170 435134
rect 412406 434898 442890 435134
rect 443126 434898 473610 435134
rect 473846 434898 504330 435134
rect 504566 434898 535050 435134
rect 535286 434898 565770 435134
rect 566006 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 89610 417454
rect 89846 417218 120330 417454
rect 120566 417218 151050 417454
rect 151286 417218 181770 417454
rect 182006 417218 212490 417454
rect 212726 417218 243210 417454
rect 243446 417218 273930 417454
rect 274166 417218 304650 417454
rect 304886 417218 335370 417454
rect 335606 417218 366090 417454
rect 366326 417218 396810 417454
rect 397046 417218 427530 417454
rect 427766 417218 458250 417454
rect 458486 417218 488970 417454
rect 489206 417218 519690 417454
rect 519926 417218 550410 417454
rect 550646 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 89610 417134
rect 89846 416898 120330 417134
rect 120566 416898 151050 417134
rect 151286 416898 181770 417134
rect 182006 416898 212490 417134
rect 212726 416898 243210 417134
rect 243446 416898 273930 417134
rect 274166 416898 304650 417134
rect 304886 416898 335370 417134
rect 335606 416898 366090 417134
rect 366326 416898 396810 417134
rect 397046 416898 427530 417134
rect 427766 416898 458250 417134
rect 458486 416898 488970 417134
rect 489206 416898 519690 417134
rect 519926 416898 550410 417134
rect 550646 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 74250 399454
rect 74486 399218 104970 399454
rect 105206 399218 135690 399454
rect 135926 399218 166410 399454
rect 166646 399218 197130 399454
rect 197366 399218 227850 399454
rect 228086 399218 258570 399454
rect 258806 399218 289290 399454
rect 289526 399218 320010 399454
rect 320246 399218 350730 399454
rect 350966 399218 381450 399454
rect 381686 399218 412170 399454
rect 412406 399218 442890 399454
rect 443126 399218 473610 399454
rect 473846 399218 504330 399454
rect 504566 399218 535050 399454
rect 535286 399218 565770 399454
rect 566006 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 74250 399134
rect 74486 398898 104970 399134
rect 105206 398898 135690 399134
rect 135926 398898 166410 399134
rect 166646 398898 197130 399134
rect 197366 398898 227850 399134
rect 228086 398898 258570 399134
rect 258806 398898 289290 399134
rect 289526 398898 320010 399134
rect 320246 398898 350730 399134
rect 350966 398898 381450 399134
rect 381686 398898 412170 399134
rect 412406 398898 442890 399134
rect 443126 398898 473610 399134
rect 473846 398898 504330 399134
rect 504566 398898 535050 399134
rect 535286 398898 565770 399134
rect 566006 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 89610 381454
rect 89846 381218 120330 381454
rect 120566 381218 151050 381454
rect 151286 381218 181770 381454
rect 182006 381218 212490 381454
rect 212726 381218 243210 381454
rect 243446 381218 273930 381454
rect 274166 381218 304650 381454
rect 304886 381218 335370 381454
rect 335606 381218 366090 381454
rect 366326 381218 396810 381454
rect 397046 381218 427530 381454
rect 427766 381218 458250 381454
rect 458486 381218 488970 381454
rect 489206 381218 519690 381454
rect 519926 381218 550410 381454
rect 550646 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 89610 381134
rect 89846 380898 120330 381134
rect 120566 380898 151050 381134
rect 151286 380898 181770 381134
rect 182006 380898 212490 381134
rect 212726 380898 243210 381134
rect 243446 380898 273930 381134
rect 274166 380898 304650 381134
rect 304886 380898 335370 381134
rect 335606 380898 366090 381134
rect 366326 380898 396810 381134
rect 397046 380898 427530 381134
rect 427766 380898 458250 381134
rect 458486 380898 488970 381134
rect 489206 380898 519690 381134
rect 519926 380898 550410 381134
rect 550646 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 135690 363454
rect 135926 363218 166410 363454
rect 166646 363218 197130 363454
rect 197366 363218 227850 363454
rect 228086 363218 258570 363454
rect 258806 363218 289290 363454
rect 289526 363218 320010 363454
rect 320246 363218 350730 363454
rect 350966 363218 381450 363454
rect 381686 363218 412170 363454
rect 412406 363218 442890 363454
rect 443126 363218 473610 363454
rect 473846 363218 504330 363454
rect 504566 363218 535050 363454
rect 535286 363218 565770 363454
rect 566006 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 135690 363134
rect 135926 362898 166410 363134
rect 166646 362898 197130 363134
rect 197366 362898 227850 363134
rect 228086 362898 258570 363134
rect 258806 362898 289290 363134
rect 289526 362898 320010 363134
rect 320246 362898 350730 363134
rect 350966 362898 381450 363134
rect 381686 362898 412170 363134
rect 412406 362898 442890 363134
rect 443126 362898 473610 363134
rect 473846 362898 504330 363134
rect 504566 362898 535050 363134
rect 535286 362898 565770 363134
rect 566006 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 120330 345454
rect 120566 345218 151050 345454
rect 151286 345218 181770 345454
rect 182006 345218 212490 345454
rect 212726 345218 243210 345454
rect 243446 345218 273930 345454
rect 274166 345218 304650 345454
rect 304886 345218 335370 345454
rect 335606 345218 366090 345454
rect 366326 345218 396810 345454
rect 397046 345218 427530 345454
rect 427766 345218 458250 345454
rect 458486 345218 488970 345454
rect 489206 345218 519690 345454
rect 519926 345218 550410 345454
rect 550646 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 120330 345134
rect 120566 344898 151050 345134
rect 151286 344898 181770 345134
rect 182006 344898 212490 345134
rect 212726 344898 243210 345134
rect 243446 344898 273930 345134
rect 274166 344898 304650 345134
rect 304886 344898 335370 345134
rect 335606 344898 366090 345134
rect 366326 344898 396810 345134
rect 397046 344898 427530 345134
rect 427766 344898 458250 345134
rect 458486 344898 488970 345134
rect 489206 344898 519690 345134
rect 519926 344898 550410 345134
rect 550646 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 74250 327454
rect 74486 327218 104970 327454
rect 105206 327218 135690 327454
rect 135926 327218 166410 327454
rect 166646 327218 197130 327454
rect 197366 327218 227850 327454
rect 228086 327218 258570 327454
rect 258806 327218 289290 327454
rect 289526 327218 320010 327454
rect 320246 327218 350730 327454
rect 350966 327218 381450 327454
rect 381686 327218 412170 327454
rect 412406 327218 442890 327454
rect 443126 327218 473610 327454
rect 473846 327218 504330 327454
rect 504566 327218 535050 327454
rect 535286 327218 565770 327454
rect 566006 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 74250 327134
rect 74486 326898 104970 327134
rect 105206 326898 135690 327134
rect 135926 326898 166410 327134
rect 166646 326898 197130 327134
rect 197366 326898 227850 327134
rect 228086 326898 258570 327134
rect 258806 326898 289290 327134
rect 289526 326898 320010 327134
rect 320246 326898 350730 327134
rect 350966 326898 381450 327134
rect 381686 326898 412170 327134
rect 412406 326898 442890 327134
rect 443126 326898 473610 327134
rect 473846 326898 504330 327134
rect 504566 326898 535050 327134
rect 535286 326898 565770 327134
rect 566006 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 89610 309454
rect 89846 309218 120330 309454
rect 120566 309218 151050 309454
rect 151286 309218 181770 309454
rect 182006 309218 212490 309454
rect 212726 309218 243210 309454
rect 243446 309218 273930 309454
rect 274166 309218 304650 309454
rect 304886 309218 335370 309454
rect 335606 309218 366090 309454
rect 366326 309218 396810 309454
rect 397046 309218 427530 309454
rect 427766 309218 458250 309454
rect 458486 309218 488970 309454
rect 489206 309218 519690 309454
rect 519926 309218 550410 309454
rect 550646 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 89610 309134
rect 89846 308898 120330 309134
rect 120566 308898 151050 309134
rect 151286 308898 181770 309134
rect 182006 308898 212490 309134
rect 212726 308898 243210 309134
rect 243446 308898 273930 309134
rect 274166 308898 304650 309134
rect 304886 308898 335370 309134
rect 335606 308898 366090 309134
rect 366326 308898 396810 309134
rect 397046 308898 427530 309134
rect 427766 308898 458250 309134
rect 458486 308898 488970 309134
rect 489206 308898 519690 309134
rect 519926 308898 550410 309134
rect 550646 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 74250 291454
rect 74486 291218 104970 291454
rect 105206 291218 135690 291454
rect 135926 291218 166410 291454
rect 166646 291218 197130 291454
rect 197366 291218 227850 291454
rect 228086 291218 258570 291454
rect 258806 291218 289290 291454
rect 289526 291218 320010 291454
rect 320246 291218 350730 291454
rect 350966 291218 381450 291454
rect 381686 291218 412170 291454
rect 412406 291218 442890 291454
rect 443126 291218 473610 291454
rect 473846 291218 504330 291454
rect 504566 291218 535050 291454
rect 535286 291218 565770 291454
rect 566006 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 74250 291134
rect 74486 290898 104970 291134
rect 105206 290898 135690 291134
rect 135926 290898 166410 291134
rect 166646 290898 197130 291134
rect 197366 290898 227850 291134
rect 228086 290898 258570 291134
rect 258806 290898 289290 291134
rect 289526 290898 320010 291134
rect 320246 290898 350730 291134
rect 350966 290898 381450 291134
rect 381686 290898 412170 291134
rect 412406 290898 442890 291134
rect 443126 290898 473610 291134
rect 473846 290898 504330 291134
rect 504566 290898 535050 291134
rect 535286 290898 565770 291134
rect 566006 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 120330 273454
rect 120566 273218 151050 273454
rect 151286 273218 181770 273454
rect 182006 273218 212490 273454
rect 212726 273218 243210 273454
rect 243446 273218 273930 273454
rect 274166 273218 304650 273454
rect 304886 273218 335370 273454
rect 335606 273218 366090 273454
rect 366326 273218 396810 273454
rect 397046 273218 427530 273454
rect 427766 273218 458250 273454
rect 458486 273218 488970 273454
rect 489206 273218 519690 273454
rect 519926 273218 550410 273454
rect 550646 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 120330 273134
rect 120566 272898 151050 273134
rect 151286 272898 181770 273134
rect 182006 272898 212490 273134
rect 212726 272898 243210 273134
rect 243446 272898 273930 273134
rect 274166 272898 304650 273134
rect 304886 272898 335370 273134
rect 335606 272898 366090 273134
rect 366326 272898 396810 273134
rect 397046 272898 427530 273134
rect 427766 272898 458250 273134
rect 458486 272898 488970 273134
rect 489206 272898 519690 273134
rect 519926 272898 550410 273134
rect 550646 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 135690 255454
rect 135926 255218 166410 255454
rect 166646 255218 197130 255454
rect 197366 255218 227850 255454
rect 228086 255218 258570 255454
rect 258806 255218 289290 255454
rect 289526 255218 320010 255454
rect 320246 255218 350730 255454
rect 350966 255218 381450 255454
rect 381686 255218 412170 255454
rect 412406 255218 442890 255454
rect 443126 255218 473610 255454
rect 473846 255218 504330 255454
rect 504566 255218 535050 255454
rect 535286 255218 565770 255454
rect 566006 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 135690 255134
rect 135926 254898 166410 255134
rect 166646 254898 197130 255134
rect 197366 254898 227850 255134
rect 228086 254898 258570 255134
rect 258806 254898 289290 255134
rect 289526 254898 320010 255134
rect 320246 254898 350730 255134
rect 350966 254898 381450 255134
rect 381686 254898 412170 255134
rect 412406 254898 442890 255134
rect 443126 254898 473610 255134
rect 473846 254898 504330 255134
rect 504566 254898 535050 255134
rect 535286 254898 565770 255134
rect 566006 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 89610 237454
rect 89846 237218 120330 237454
rect 120566 237218 151050 237454
rect 151286 237218 181770 237454
rect 182006 237218 212490 237454
rect 212726 237218 243210 237454
rect 243446 237218 273930 237454
rect 274166 237218 304650 237454
rect 304886 237218 335370 237454
rect 335606 237218 366090 237454
rect 366326 237218 396810 237454
rect 397046 237218 427530 237454
rect 427766 237218 458250 237454
rect 458486 237218 488970 237454
rect 489206 237218 519690 237454
rect 519926 237218 550410 237454
rect 550646 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 89610 237134
rect 89846 236898 120330 237134
rect 120566 236898 151050 237134
rect 151286 236898 181770 237134
rect 182006 236898 212490 237134
rect 212726 236898 243210 237134
rect 243446 236898 273930 237134
rect 274166 236898 304650 237134
rect 304886 236898 335370 237134
rect 335606 236898 366090 237134
rect 366326 236898 396810 237134
rect 397046 236898 427530 237134
rect 427766 236898 458250 237134
rect 458486 236898 488970 237134
rect 489206 236898 519690 237134
rect 519926 236898 550410 237134
rect 550646 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 74250 219454
rect 74486 219218 104970 219454
rect 105206 219218 135690 219454
rect 135926 219218 166410 219454
rect 166646 219218 197130 219454
rect 197366 219218 227850 219454
rect 228086 219218 258570 219454
rect 258806 219218 289290 219454
rect 289526 219218 320010 219454
rect 320246 219218 350730 219454
rect 350966 219218 381450 219454
rect 381686 219218 412170 219454
rect 412406 219218 442890 219454
rect 443126 219218 473610 219454
rect 473846 219218 504330 219454
rect 504566 219218 535050 219454
rect 535286 219218 565770 219454
rect 566006 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 74250 219134
rect 74486 218898 104970 219134
rect 105206 218898 135690 219134
rect 135926 218898 166410 219134
rect 166646 218898 197130 219134
rect 197366 218898 227850 219134
rect 228086 218898 258570 219134
rect 258806 218898 289290 219134
rect 289526 218898 320010 219134
rect 320246 218898 350730 219134
rect 350966 218898 381450 219134
rect 381686 218898 412170 219134
rect 412406 218898 442890 219134
rect 443126 218898 473610 219134
rect 473846 218898 504330 219134
rect 504566 218898 535050 219134
rect 535286 218898 565770 219134
rect 566006 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 89610 201454
rect 89846 201218 120330 201454
rect 120566 201218 151050 201454
rect 151286 201218 181770 201454
rect 182006 201218 212490 201454
rect 212726 201218 243210 201454
rect 243446 201218 273930 201454
rect 274166 201218 304650 201454
rect 304886 201218 335370 201454
rect 335606 201218 366090 201454
rect 366326 201218 396810 201454
rect 397046 201218 427530 201454
rect 427766 201218 458250 201454
rect 458486 201218 488970 201454
rect 489206 201218 519690 201454
rect 519926 201218 550410 201454
rect 550646 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 89610 201134
rect 89846 200898 120330 201134
rect 120566 200898 151050 201134
rect 151286 200898 181770 201134
rect 182006 200898 212490 201134
rect 212726 200898 243210 201134
rect 243446 200898 273930 201134
rect 274166 200898 304650 201134
rect 304886 200898 335370 201134
rect 335606 200898 366090 201134
rect 366326 200898 396810 201134
rect 397046 200898 427530 201134
rect 427766 200898 458250 201134
rect 458486 200898 488970 201134
rect 489206 200898 519690 201134
rect 519926 200898 550410 201134
rect 550646 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 74250 183454
rect 74486 183218 104970 183454
rect 105206 183218 135690 183454
rect 135926 183218 166410 183454
rect 166646 183218 197130 183454
rect 197366 183218 227850 183454
rect 228086 183218 258570 183454
rect 258806 183218 289290 183454
rect 289526 183218 320010 183454
rect 320246 183218 350730 183454
rect 350966 183218 381450 183454
rect 381686 183218 412170 183454
rect 412406 183218 442890 183454
rect 443126 183218 473610 183454
rect 473846 183218 504330 183454
rect 504566 183218 535050 183454
rect 535286 183218 565770 183454
rect 566006 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 74250 183134
rect 74486 182898 104970 183134
rect 105206 182898 135690 183134
rect 135926 182898 166410 183134
rect 166646 182898 197130 183134
rect 197366 182898 227850 183134
rect 228086 182898 258570 183134
rect 258806 182898 289290 183134
rect 289526 182898 320010 183134
rect 320246 182898 350730 183134
rect 350966 182898 381450 183134
rect 381686 182898 412170 183134
rect 412406 182898 442890 183134
rect 443126 182898 473610 183134
rect 473846 182898 504330 183134
rect 504566 182898 535050 183134
rect 535286 182898 565770 183134
rect 566006 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 89610 165454
rect 89846 165218 120330 165454
rect 120566 165218 151050 165454
rect 151286 165218 181770 165454
rect 182006 165218 212490 165454
rect 212726 165218 243210 165454
rect 243446 165218 273930 165454
rect 274166 165218 304650 165454
rect 304886 165218 335370 165454
rect 335606 165218 366090 165454
rect 366326 165218 396810 165454
rect 397046 165218 427530 165454
rect 427766 165218 458250 165454
rect 458486 165218 488970 165454
rect 489206 165218 519690 165454
rect 519926 165218 550410 165454
rect 550646 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 89610 165134
rect 89846 164898 120330 165134
rect 120566 164898 151050 165134
rect 151286 164898 181770 165134
rect 182006 164898 212490 165134
rect 212726 164898 243210 165134
rect 243446 164898 273930 165134
rect 274166 164898 304650 165134
rect 304886 164898 335370 165134
rect 335606 164898 366090 165134
rect 366326 164898 396810 165134
rect 397046 164898 427530 165134
rect 427766 164898 458250 165134
rect 458486 164898 488970 165134
rect 489206 164898 519690 165134
rect 519926 164898 550410 165134
rect 550646 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 74250 147454
rect 74486 147218 104970 147454
rect 105206 147218 135690 147454
rect 135926 147218 166410 147454
rect 166646 147218 197130 147454
rect 197366 147218 227850 147454
rect 228086 147218 258570 147454
rect 258806 147218 289290 147454
rect 289526 147218 320010 147454
rect 320246 147218 350730 147454
rect 350966 147218 381450 147454
rect 381686 147218 412170 147454
rect 412406 147218 442890 147454
rect 443126 147218 473610 147454
rect 473846 147218 504330 147454
rect 504566 147218 535050 147454
rect 535286 147218 565770 147454
rect 566006 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 74250 147134
rect 74486 146898 104970 147134
rect 105206 146898 135690 147134
rect 135926 146898 166410 147134
rect 166646 146898 197130 147134
rect 197366 146898 227850 147134
rect 228086 146898 258570 147134
rect 258806 146898 289290 147134
rect 289526 146898 320010 147134
rect 320246 146898 350730 147134
rect 350966 146898 381450 147134
rect 381686 146898 412170 147134
rect 412406 146898 442890 147134
rect 443126 146898 473610 147134
rect 473846 146898 504330 147134
rect 504566 146898 535050 147134
rect 535286 146898 565770 147134
rect 566006 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 89610 129454
rect 89846 129218 120330 129454
rect 120566 129218 151050 129454
rect 151286 129218 181770 129454
rect 182006 129218 212490 129454
rect 212726 129218 243210 129454
rect 243446 129218 273930 129454
rect 274166 129218 304650 129454
rect 304886 129218 335370 129454
rect 335606 129218 366090 129454
rect 366326 129218 396810 129454
rect 397046 129218 427530 129454
rect 427766 129218 458250 129454
rect 458486 129218 488970 129454
rect 489206 129218 519690 129454
rect 519926 129218 550410 129454
rect 550646 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 89610 129134
rect 89846 128898 120330 129134
rect 120566 128898 151050 129134
rect 151286 128898 181770 129134
rect 182006 128898 212490 129134
rect 212726 128898 243210 129134
rect 243446 128898 273930 129134
rect 274166 128898 304650 129134
rect 304886 128898 335370 129134
rect 335606 128898 366090 129134
rect 366326 128898 396810 129134
rect 397046 128898 427530 129134
rect 427766 128898 458250 129134
rect 458486 128898 488970 129134
rect 489206 128898 519690 129134
rect 519926 128898 550410 129134
rect 550646 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 74250 111454
rect 74486 111218 104970 111454
rect 105206 111218 135690 111454
rect 135926 111218 166410 111454
rect 166646 111218 197130 111454
rect 197366 111218 227850 111454
rect 228086 111218 258570 111454
rect 258806 111218 289290 111454
rect 289526 111218 320010 111454
rect 320246 111218 350730 111454
rect 350966 111218 381450 111454
rect 381686 111218 412170 111454
rect 412406 111218 442890 111454
rect 443126 111218 473610 111454
rect 473846 111218 504330 111454
rect 504566 111218 535050 111454
rect 535286 111218 565770 111454
rect 566006 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 74250 111134
rect 74486 110898 104970 111134
rect 105206 110898 135690 111134
rect 135926 110898 166410 111134
rect 166646 110898 197130 111134
rect 197366 110898 227850 111134
rect 228086 110898 258570 111134
rect 258806 110898 289290 111134
rect 289526 110898 320010 111134
rect 320246 110898 350730 111134
rect 350966 110898 381450 111134
rect 381686 110898 412170 111134
rect 412406 110898 442890 111134
rect 443126 110898 473610 111134
rect 473846 110898 504330 111134
rect 504566 110898 535050 111134
rect 535286 110898 565770 111134
rect 566006 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 89610 93454
rect 89846 93218 120330 93454
rect 120566 93218 151050 93454
rect 151286 93218 181770 93454
rect 182006 93218 212490 93454
rect 212726 93218 243210 93454
rect 243446 93218 273930 93454
rect 274166 93218 304650 93454
rect 304886 93218 335370 93454
rect 335606 93218 366090 93454
rect 366326 93218 396810 93454
rect 397046 93218 427530 93454
rect 427766 93218 458250 93454
rect 458486 93218 488970 93454
rect 489206 93218 519690 93454
rect 519926 93218 550410 93454
rect 550646 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 89610 93134
rect 89846 92898 120330 93134
rect 120566 92898 151050 93134
rect 151286 92898 181770 93134
rect 182006 92898 212490 93134
rect 212726 92898 243210 93134
rect 243446 92898 273930 93134
rect 274166 92898 304650 93134
rect 304886 92898 335370 93134
rect 335606 92898 366090 93134
rect 366326 92898 396810 93134
rect 397046 92898 427530 93134
rect 427766 92898 458250 93134
rect 458486 92898 488970 93134
rect 489206 92898 519690 93134
rect 519926 92898 550410 93134
rect 550646 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 74250 75454
rect 74486 75218 104970 75454
rect 105206 75218 135690 75454
rect 135926 75218 166410 75454
rect 166646 75218 197130 75454
rect 197366 75218 227850 75454
rect 228086 75218 258570 75454
rect 258806 75218 289290 75454
rect 289526 75218 320010 75454
rect 320246 75218 350730 75454
rect 350966 75218 381450 75454
rect 381686 75218 412170 75454
rect 412406 75218 442890 75454
rect 443126 75218 473610 75454
rect 473846 75218 504330 75454
rect 504566 75218 535050 75454
rect 535286 75218 565770 75454
rect 566006 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 74250 75134
rect 74486 74898 104970 75134
rect 105206 74898 135690 75134
rect 135926 74898 166410 75134
rect 166646 74898 197130 75134
rect 197366 74898 227850 75134
rect 228086 74898 258570 75134
rect 258806 74898 289290 75134
rect 289526 74898 320010 75134
rect 320246 74898 350730 75134
rect 350966 74898 381450 75134
rect 381686 74898 412170 75134
rect 412406 74898 442890 75134
rect 443126 74898 473610 75134
rect 473846 74898 504330 75134
rect 504566 74898 535050 75134
rect 535286 74898 565770 75134
rect 566006 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use both  both
timestamp 1641005295
transform 1 0 70000 0 1 68000
box -10 0 500000 500000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 66000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 570000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 570000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 570000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 570000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 570000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 570000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 570000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 570000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 570000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 570000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 570000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 570000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 570000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 570000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 66000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 570000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 570000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 570000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 570000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 570000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 570000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 570000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 570000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 570000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 570000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 570000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 570000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 570000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 570000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 66000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 570000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 570000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 570000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 570000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 570000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 570000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 570000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 570000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 570000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 570000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 570000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 570000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 570000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 570000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 66000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 570000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 570000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 570000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 570000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 570000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 570000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 570000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 570000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 570000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 570000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 570000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 570000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 570000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 570000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 66000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 570000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 570000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 570000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 570000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 570000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 570000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 570000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 570000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 570000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 570000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 570000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 570000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 570000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 570000 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 66000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 570000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 570000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 570000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 570000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 570000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 570000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 570000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 570000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 570000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 570000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 570000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 570000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 570000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 570000 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 66000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 570000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 570000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 570000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 570000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 570000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 570000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 570000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 570000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 570000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 570000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 570000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 570000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 570000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 570000 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 66000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 570000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 570000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 570000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 570000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 570000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 570000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 570000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 570000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 570000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 570000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 570000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 570000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 570000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 570000 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
