VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO both
  CLASS BLOCK ;
  FOREIGN both ;
  ORIGIN 0.000 0.000 ;
  SIZE 289.020 BY 299.740 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 0.000 96.190 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.100 4.000 206.300 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 295.740 8.790 299.740 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 273.100 289.020 274.300 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.990 295.740 11.550 299.740 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 295.740 104.470 299.740 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 0.000 152.310 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.790 295.740 117.350 299.740 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 295.740 269.150 299.740 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.190 0.000 89.750 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 269.020 289.020 270.220 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.540 4.000 279.740 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 295.740 151.390 299.740 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 0.000 139.430 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.430 295.740 17.990 299.740 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 39.180 289.020 40.380 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 213.260 289.020 214.460 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.300 4.000 165.500 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 295.740 82.390 299.740 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 0.000 34.550 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.420 4.000 188.620 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 295.740 169.790 299.740 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 0.000 186.350 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 254.060 289.020 255.260 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.900 4.000 179.100 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.910 0.000 12.470 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.060 4.000 119.260 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 79.980 289.020 81.180 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 295.740 76.870 299.740 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 295.740 23.510 299.740 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.270 0.000 111.830 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 295.740 215.790 299.740 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.630 295.740 188.190 299.740 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 295.740 73.190 299.740 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 290.780 289.020 291.980 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.270 295.740 249.830 299.740 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.780 4.000 155.980 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 295.740 228.670 299.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 222.780 289.020 223.980 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.220 4.000 229.420 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 135.740 289.020 136.940 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 0.000 30.870 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.310 0.000 260.870 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 295.740 61.230 299.740 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.860 4.000 160.060 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 71.820 289.020 73.020 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.220 4.000 59.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 295.740 138.510 299.740 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 295.740 107.230 299.740 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 0.000 114.590 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.820 4.000 5.020 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 0.000 83.310 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 0.000 247.990 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.980 4.000 183.180 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 162.940 289.020 164.140 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.230 0.000 284.790 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 0.000 220.390 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.780 4.000 87.980 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 181.980 289.020 183.180 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 0.000 68.590 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.350 295.740 110.910 299.740 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 295.740 247.070 299.740 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 186.060 289.020 187.260 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 0.000 136.670 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 0.000 288.470 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.830 0.000 59.390 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 66.380 289.020 67.580 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 295.740 135.750 299.740 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.900 4.000 247.100 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.500 4.000 22.700 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 295.740 144.950 299.740 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.510 0.000 270.070 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 149.340 289.020 150.540 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 295.740 86.070 299.740 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 0.000 223.150 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.620 4.000 283.820 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 158.860 289.020 160.060 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 296.220 289.020 297.420 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.710 295.740 141.270 299.740 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 218.700 289.020 219.900 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 295.740 231.430 299.740 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 295.740 281.110 299.740 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.950 295.740 92.510 299.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 58.220 289.020 59.420 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 295.740 200.150 299.740 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 295.740 283.870 299.740 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.700 4.000 151.900 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.870 0.000 254.430 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 62.300 289.020 63.500 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 0.000 204.750 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 295.740 48.350 299.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.350 0.000 179.910 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 0.000 21.670 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 295.740 20.750 299.740 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 108.540 289.020 109.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 0.000 62.150 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230 0.000 238.790 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.500 4.000 192.700 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.060 4.000 289.260 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 295.740 166.110 299.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.710 295.740 210.270 299.740 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 0.000 46.510 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 245.900 289.020 247.100 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.990 295.740 172.550 299.740 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.910 0.000 173.470 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 0.000 195.550 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.590 0.000 108.150 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 295.740 194.630 299.740 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 167.020 289.020 168.220 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 44.620 289.020 45.820 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 295.740 98.030 299.740 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 295.740 29.950 299.740 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 295.740 45.590 299.740 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.980 4.000 115.180 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.260 4.000 78.460 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.270 0.000 272.830 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 203.740 289.020 204.940 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 0.000 15.230 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 0.000 98.950 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 295.740 274.670 299.740 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 295.740 113.670 299.740 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 0.000 225.910 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 295.740 88.830 299.740 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.020 4.000 32.220 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 89.500 289.020 90.700 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 282.620 289.020 283.820 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.220 4.000 297.420 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.300 4.000 233.500 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.510 0.000 201.070 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.990 0.000 241.550 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 145.260 289.020 146.460 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.590 295.740 154.150 299.740 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.470 0.000 282.030 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.070 0.000 263.630 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 295.740 156.910 299.740 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 16.060 289.020 17.260 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.060 4.000 51.260 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 21.500 289.020 22.700 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.420 4.000 256.620 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.070 295.740 33.630 299.740 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 0.000 43.750 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 0.000 155.070 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 295.740 237.870 299.740 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 295.740 120.110 299.740 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 176.540 289.020 177.740 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 232.300 289.020 233.500 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.150 295.740 147.710 299.740 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.860 4.000 92.060 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 295.740 39.150 299.740 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 295.740 79.630 299.740 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.020 4.000 270.220 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.620 4.000 215.820 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 153.420 289.020 154.620 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 172.460 289.020 173.660 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.470 295.740 259.030 299.740 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 116.700 289.020 117.900 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.070 0.000 102.630 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 295.740 14.310 299.740 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 295.740 224.990 299.740 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.580 4.000 128.780 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.830 0.000 105.390 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.390 0.000 213.950 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 195.580 289.020 196.780 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 0.000 6.030 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 0.000 40.070 4.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.670 295.740 176.230 299.740 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.470 0.000 167.030 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 0.000 80.550 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 0.000 157.830 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 35.100 289.020 36.300 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.140 4.000 293.340 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.710 0.000 164.270 4.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 295.740 213.030 299.740 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 0.000 211.190 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 85.420 289.020 86.620 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.990 295.740 287.550 299.740 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 48.700 289.020 49.900 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.180 4.000 210.380 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 240.460 289.020 241.660 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 0.000 236.030 4.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.150 295.740 262.710 299.740 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 0.000 198.310 4.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.870 295.740 185.430 299.740 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 0.000 28.110 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.550 295.740 5.110 299.740 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 0.000 121.030 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.230 295.740 54.790 299.740 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 0.000 55.710 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.950 0.000 207.510 4.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 295.740 190.950 299.740 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 263.580 289.020 264.780 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.150 295.740 101.710 299.740 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 295.740 58.470 299.740 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 295.740 197.390 299.740 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 0.000 257.190 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.030 295.740 160.590 299.740 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 11.980 289.020 13.180 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 295.740 265.470 299.740 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 295.740 219.470 299.740 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 295.740 67.670 299.740 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.820 4.000 175.020 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.430 295.740 63.990 299.740 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 139.820 289.020 141.020 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 122.140 289.020 123.340 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 99.020 289.020 100.220 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 7.900 289.020 9.100 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.150 0.000 216.710 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.950 295.740 253.510 299.740 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 259.500 289.020 260.700 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.910 0.000 127.470 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 0.000 182.670 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.030 0.000 275.590 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 295.740 129.310 299.740 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 0.000 123.790 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.870 0.000 24.430 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 295.740 178.990 299.740 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 103.100 289.020 104.300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 226.860 289.020 228.060 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 0.000 86.990 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790 295.740 278.350 299.740 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 52.780 289.020 53.980 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.420 4.000 18.620 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.150 0.000 170.710 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 0.000 71.350 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030 0.000 229.590 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 2.460 289.020 3.660 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.790 295.740 163.350 299.740 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.660 4.000 64.860 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 295.740 36.390 299.740 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 295.740 52.030 299.740 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 295.740 42.830 299.740 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.380 4.000 101.580 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 94.940 289.020 96.140 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 0.000 132.990 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.070 295.740 240.630 299.740 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 286.700 289.020 287.900 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 295.740 95.270 299.740 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 277.180 289.020 278.380 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.460 4.000 275.660 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 190.140 289.020 191.340 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.350 295.740 271.910 299.740 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.510 295.740 132.070 299.740 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 0.000 74.110 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 131.660 289.020 132.860 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.310 0.000 191.870 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 25.580 289.020 26.780 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.820 4.000 243.020 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 0.000 245.230 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.750 0.000 37.310 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.710 0.000 118.270 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 75.900 289.020 77.100 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 295.740 256.270 299.740 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 236.380 289.020 237.580 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 0.000 250.750 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 126.220 289.020 127.420 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 0.000 3.270 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 249.980 289.020 251.180 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 295.740 244.310 299.740 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 0.000 266.390 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 295.740 235.110 299.740 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.660 4.000 132.860 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.260 4.000 146.460 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 0.000 161.510 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.550 0.000 189.110 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.580 4.000 196.780 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 295.740 122.870 299.740 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.180 4.000 142.380 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 295.740 181.750 299.740 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 295.740 126.550 299.740 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.670 0.000 130.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.670 295.740 222.230 299.740 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 29.660 289.020 30.860 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.340 4.000 252.540 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 209.180 289.020 210.380 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.390 0.000 52.950 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 0.000 93.430 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 0.000 145.870 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 199.660 289.020 200.860 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 0.000 148.630 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 295.740 206.590 299.740 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 295.740 203.830 299.740 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.630 295.740 27.190 299.740 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.870 295.740 70.430 299.740 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 0.000 177.150 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 295.740 2.350 299.740 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.020 112.620 289.020 113.820 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 3.825 0.085 288.735 296.735 ;
      LAYER met1 ;
        RECT 0.070 0.040 288.810 296.780 ;
      LAYER met2 ;
        RECT 0.100 295.460 1.510 297.005 ;
        RECT 2.630 295.460 4.270 297.005 ;
        RECT 5.390 295.460 7.950 297.005 ;
        RECT 9.070 295.460 10.710 297.005 ;
        RECT 11.830 295.460 13.470 297.005 ;
        RECT 14.590 295.460 17.150 297.005 ;
        RECT 18.270 295.460 19.910 297.005 ;
        RECT 21.030 295.460 22.670 297.005 ;
        RECT 23.790 295.460 26.350 297.005 ;
        RECT 27.470 295.460 29.110 297.005 ;
        RECT 30.230 295.460 32.790 297.005 ;
        RECT 33.910 295.460 35.550 297.005 ;
        RECT 36.670 295.460 38.310 297.005 ;
        RECT 39.430 295.460 41.990 297.005 ;
        RECT 43.110 295.460 44.750 297.005 ;
        RECT 45.870 295.460 47.510 297.005 ;
        RECT 48.630 295.460 51.190 297.005 ;
        RECT 52.310 295.460 53.950 297.005 ;
        RECT 55.070 295.460 57.630 297.005 ;
        RECT 58.750 295.460 60.390 297.005 ;
        RECT 61.510 295.460 63.150 297.005 ;
        RECT 64.270 295.460 66.830 297.005 ;
        RECT 67.950 295.460 69.590 297.005 ;
        RECT 70.710 295.460 72.350 297.005 ;
        RECT 73.470 295.460 76.030 297.005 ;
        RECT 77.150 295.460 78.790 297.005 ;
        RECT 79.910 295.460 81.550 297.005 ;
        RECT 82.670 295.460 85.230 297.005 ;
        RECT 86.350 295.460 87.990 297.005 ;
        RECT 89.110 295.460 91.670 297.005 ;
        RECT 92.790 295.460 94.430 297.005 ;
        RECT 95.550 295.460 97.190 297.005 ;
        RECT 98.310 295.460 100.870 297.005 ;
        RECT 101.990 295.460 103.630 297.005 ;
        RECT 104.750 295.460 106.390 297.005 ;
        RECT 107.510 295.460 110.070 297.005 ;
        RECT 111.190 295.460 112.830 297.005 ;
        RECT 113.950 295.460 116.510 297.005 ;
        RECT 117.630 295.460 119.270 297.005 ;
        RECT 120.390 295.460 122.030 297.005 ;
        RECT 123.150 295.460 125.710 297.005 ;
        RECT 126.830 295.460 128.470 297.005 ;
        RECT 129.590 295.460 131.230 297.005 ;
        RECT 132.350 295.460 134.910 297.005 ;
        RECT 136.030 295.460 137.670 297.005 ;
        RECT 138.790 295.460 140.430 297.005 ;
        RECT 141.550 295.460 144.110 297.005 ;
        RECT 145.230 295.460 146.870 297.005 ;
        RECT 147.990 295.460 150.550 297.005 ;
        RECT 151.670 295.460 153.310 297.005 ;
        RECT 154.430 295.460 156.070 297.005 ;
        RECT 157.190 295.460 159.750 297.005 ;
        RECT 160.870 295.460 162.510 297.005 ;
        RECT 163.630 295.460 165.270 297.005 ;
        RECT 166.390 295.460 168.950 297.005 ;
        RECT 170.070 295.460 171.710 297.005 ;
        RECT 172.830 295.460 175.390 297.005 ;
        RECT 176.510 295.460 178.150 297.005 ;
        RECT 179.270 295.460 180.910 297.005 ;
        RECT 182.030 295.460 184.590 297.005 ;
        RECT 185.710 295.460 187.350 297.005 ;
        RECT 188.470 295.460 190.110 297.005 ;
        RECT 191.230 295.460 193.790 297.005 ;
        RECT 194.910 295.460 196.550 297.005 ;
        RECT 197.670 295.460 199.310 297.005 ;
        RECT 200.430 295.460 202.990 297.005 ;
        RECT 204.110 295.460 205.750 297.005 ;
        RECT 206.870 295.460 209.430 297.005 ;
        RECT 210.550 295.460 212.190 297.005 ;
        RECT 213.310 295.460 214.950 297.005 ;
        RECT 216.070 295.460 218.630 297.005 ;
        RECT 219.750 295.460 221.390 297.005 ;
        RECT 222.510 295.460 224.150 297.005 ;
        RECT 225.270 295.460 227.830 297.005 ;
        RECT 228.950 295.460 230.590 297.005 ;
        RECT 231.710 295.460 234.270 297.005 ;
        RECT 235.390 295.460 237.030 297.005 ;
        RECT 238.150 295.460 239.790 297.005 ;
        RECT 240.910 295.460 243.470 297.005 ;
        RECT 244.590 295.460 246.230 297.005 ;
        RECT 247.350 295.460 248.990 297.005 ;
        RECT 250.110 295.460 252.670 297.005 ;
        RECT 253.790 295.460 255.430 297.005 ;
        RECT 256.550 295.460 258.190 297.005 ;
        RECT 259.310 295.460 261.870 297.005 ;
        RECT 262.990 295.460 264.630 297.005 ;
        RECT 265.750 295.460 268.310 297.005 ;
        RECT 269.430 295.460 271.070 297.005 ;
        RECT 272.190 295.460 273.830 297.005 ;
        RECT 274.950 295.460 277.510 297.005 ;
        RECT 278.630 295.460 280.270 297.005 ;
        RECT 281.390 295.460 283.030 297.005 ;
        RECT 284.150 295.460 286.710 297.005 ;
        RECT 287.830 295.460 288.780 297.005 ;
        RECT 0.100 4.280 288.780 295.460 ;
        RECT 0.790 0.010 2.430 4.280 ;
        RECT 3.550 0.010 5.190 4.280 ;
        RECT 6.310 0.010 8.870 4.280 ;
        RECT 9.990 0.010 11.630 4.280 ;
        RECT 12.750 0.010 14.390 4.280 ;
        RECT 15.510 0.010 18.070 4.280 ;
        RECT 19.190 0.010 20.830 4.280 ;
        RECT 21.950 0.010 23.590 4.280 ;
        RECT 24.710 0.010 27.270 4.280 ;
        RECT 28.390 0.010 30.030 4.280 ;
        RECT 31.150 0.010 33.710 4.280 ;
        RECT 34.830 0.010 36.470 4.280 ;
        RECT 37.590 0.010 39.230 4.280 ;
        RECT 40.350 0.010 42.910 4.280 ;
        RECT 44.030 0.010 45.670 4.280 ;
        RECT 46.790 0.010 48.430 4.280 ;
        RECT 49.550 0.010 52.110 4.280 ;
        RECT 53.230 0.010 54.870 4.280 ;
        RECT 55.990 0.010 58.550 4.280 ;
        RECT 59.670 0.010 61.310 4.280 ;
        RECT 62.430 0.010 64.070 4.280 ;
        RECT 65.190 0.010 67.750 4.280 ;
        RECT 68.870 0.010 70.510 4.280 ;
        RECT 71.630 0.010 73.270 4.280 ;
        RECT 74.390 0.010 76.950 4.280 ;
        RECT 78.070 0.010 79.710 4.280 ;
        RECT 80.830 0.010 82.470 4.280 ;
        RECT 83.590 0.010 86.150 4.280 ;
        RECT 87.270 0.010 88.910 4.280 ;
        RECT 90.030 0.010 92.590 4.280 ;
        RECT 93.710 0.010 95.350 4.280 ;
        RECT 96.470 0.010 98.110 4.280 ;
        RECT 99.230 0.010 101.790 4.280 ;
        RECT 102.910 0.010 104.550 4.280 ;
        RECT 105.670 0.010 107.310 4.280 ;
        RECT 108.430 0.010 110.990 4.280 ;
        RECT 112.110 0.010 113.750 4.280 ;
        RECT 114.870 0.010 117.430 4.280 ;
        RECT 118.550 0.010 120.190 4.280 ;
        RECT 121.310 0.010 122.950 4.280 ;
        RECT 124.070 0.010 126.630 4.280 ;
        RECT 127.750 0.010 129.390 4.280 ;
        RECT 130.510 0.010 132.150 4.280 ;
        RECT 133.270 0.010 135.830 4.280 ;
        RECT 136.950 0.010 138.590 4.280 ;
        RECT 139.710 0.010 141.350 4.280 ;
        RECT 142.470 0.010 145.030 4.280 ;
        RECT 146.150 0.010 147.790 4.280 ;
        RECT 148.910 0.010 151.470 4.280 ;
        RECT 152.590 0.010 154.230 4.280 ;
        RECT 155.350 0.010 156.990 4.280 ;
        RECT 158.110 0.010 160.670 4.280 ;
        RECT 161.790 0.010 163.430 4.280 ;
        RECT 164.550 0.010 166.190 4.280 ;
        RECT 167.310 0.010 169.870 4.280 ;
        RECT 170.990 0.010 172.630 4.280 ;
        RECT 173.750 0.010 176.310 4.280 ;
        RECT 177.430 0.010 179.070 4.280 ;
        RECT 180.190 0.010 181.830 4.280 ;
        RECT 182.950 0.010 185.510 4.280 ;
        RECT 186.630 0.010 188.270 4.280 ;
        RECT 189.390 0.010 191.030 4.280 ;
        RECT 192.150 0.010 194.710 4.280 ;
        RECT 195.830 0.010 197.470 4.280 ;
        RECT 198.590 0.010 200.230 4.280 ;
        RECT 201.350 0.010 203.910 4.280 ;
        RECT 205.030 0.010 206.670 4.280 ;
        RECT 207.790 0.010 210.350 4.280 ;
        RECT 211.470 0.010 213.110 4.280 ;
        RECT 214.230 0.010 215.870 4.280 ;
        RECT 216.990 0.010 219.550 4.280 ;
        RECT 220.670 0.010 222.310 4.280 ;
        RECT 223.430 0.010 225.070 4.280 ;
        RECT 226.190 0.010 228.750 4.280 ;
        RECT 229.870 0.010 231.510 4.280 ;
        RECT 232.630 0.010 235.190 4.280 ;
        RECT 236.310 0.010 237.950 4.280 ;
        RECT 239.070 0.010 240.710 4.280 ;
        RECT 241.830 0.010 244.390 4.280 ;
        RECT 245.510 0.010 247.150 4.280 ;
        RECT 248.270 0.010 249.910 4.280 ;
        RECT 251.030 0.010 253.590 4.280 ;
        RECT 254.710 0.010 256.350 4.280 ;
        RECT 257.470 0.010 260.030 4.280 ;
        RECT 261.150 0.010 262.790 4.280 ;
        RECT 263.910 0.010 265.550 4.280 ;
        RECT 266.670 0.010 269.230 4.280 ;
        RECT 270.350 0.010 271.990 4.280 ;
        RECT 273.110 0.010 274.750 4.280 ;
        RECT 275.870 0.010 278.430 4.280 ;
        RECT 279.550 0.010 281.190 4.280 ;
        RECT 282.310 0.010 283.950 4.280 ;
        RECT 285.070 0.010 287.630 4.280 ;
        RECT 288.750 0.010 288.780 4.280 ;
      LAYER met3 ;
        RECT 4.400 295.820 284.620 296.985 ;
        RECT 0.270 293.740 287.435 295.820 ;
        RECT 4.400 292.380 287.435 293.740 ;
        RECT 4.400 291.740 284.620 292.380 ;
        RECT 0.270 290.380 284.620 291.740 ;
        RECT 0.270 289.660 287.435 290.380 ;
        RECT 4.400 288.300 287.435 289.660 ;
        RECT 4.400 287.660 284.620 288.300 ;
        RECT 0.270 286.300 284.620 287.660 ;
        RECT 0.270 284.220 287.435 286.300 ;
        RECT 4.400 282.220 284.620 284.220 ;
        RECT 0.270 280.140 287.435 282.220 ;
        RECT 4.400 278.780 287.435 280.140 ;
        RECT 4.400 278.140 284.620 278.780 ;
        RECT 0.270 276.780 284.620 278.140 ;
        RECT 0.270 276.060 287.435 276.780 ;
        RECT 4.400 274.700 287.435 276.060 ;
        RECT 4.400 274.060 284.620 274.700 ;
        RECT 0.270 272.700 284.620 274.060 ;
        RECT 0.270 270.620 287.435 272.700 ;
        RECT 4.400 268.620 284.620 270.620 ;
        RECT 0.270 266.540 287.435 268.620 ;
        RECT 4.400 265.180 287.435 266.540 ;
        RECT 4.400 264.540 284.620 265.180 ;
        RECT 0.270 263.180 284.620 264.540 ;
        RECT 0.270 262.460 287.435 263.180 ;
        RECT 4.400 261.100 287.435 262.460 ;
        RECT 4.400 260.460 284.620 261.100 ;
        RECT 0.270 259.100 284.620 260.460 ;
        RECT 0.270 257.020 287.435 259.100 ;
        RECT 4.400 255.660 287.435 257.020 ;
        RECT 4.400 255.020 284.620 255.660 ;
        RECT 0.270 253.660 284.620 255.020 ;
        RECT 0.270 252.940 287.435 253.660 ;
        RECT 4.400 251.580 287.435 252.940 ;
        RECT 4.400 250.940 284.620 251.580 ;
        RECT 0.270 249.580 284.620 250.940 ;
        RECT 0.270 247.500 287.435 249.580 ;
        RECT 4.400 245.500 284.620 247.500 ;
        RECT 0.270 243.420 287.435 245.500 ;
        RECT 4.400 242.060 287.435 243.420 ;
        RECT 4.400 241.420 284.620 242.060 ;
        RECT 0.270 240.060 284.620 241.420 ;
        RECT 0.270 239.340 287.435 240.060 ;
        RECT 4.400 237.980 287.435 239.340 ;
        RECT 4.400 237.340 284.620 237.980 ;
        RECT 0.270 235.980 284.620 237.340 ;
        RECT 0.270 233.900 287.435 235.980 ;
        RECT 4.400 231.900 284.620 233.900 ;
        RECT 0.270 229.820 287.435 231.900 ;
        RECT 4.400 228.460 287.435 229.820 ;
        RECT 4.400 227.820 284.620 228.460 ;
        RECT 0.270 226.460 284.620 227.820 ;
        RECT 0.270 225.740 287.435 226.460 ;
        RECT 4.400 224.380 287.435 225.740 ;
        RECT 4.400 223.740 284.620 224.380 ;
        RECT 0.270 222.380 284.620 223.740 ;
        RECT 0.270 220.300 287.435 222.380 ;
        RECT 4.400 218.300 284.620 220.300 ;
        RECT 0.270 216.220 287.435 218.300 ;
        RECT 4.400 214.860 287.435 216.220 ;
        RECT 4.400 214.220 284.620 214.860 ;
        RECT 0.270 212.860 284.620 214.220 ;
        RECT 0.270 210.780 287.435 212.860 ;
        RECT 4.400 208.780 284.620 210.780 ;
        RECT 0.270 206.700 287.435 208.780 ;
        RECT 4.400 205.340 287.435 206.700 ;
        RECT 4.400 204.700 284.620 205.340 ;
        RECT 0.270 203.340 284.620 204.700 ;
        RECT 0.270 202.620 287.435 203.340 ;
        RECT 4.400 201.260 287.435 202.620 ;
        RECT 4.400 200.620 284.620 201.260 ;
        RECT 0.270 199.260 284.620 200.620 ;
        RECT 0.270 197.180 287.435 199.260 ;
        RECT 4.400 195.180 284.620 197.180 ;
        RECT 0.270 193.100 287.435 195.180 ;
        RECT 4.400 191.740 287.435 193.100 ;
        RECT 4.400 191.100 284.620 191.740 ;
        RECT 0.270 189.740 284.620 191.100 ;
        RECT 0.270 189.020 287.435 189.740 ;
        RECT 4.400 187.660 287.435 189.020 ;
        RECT 4.400 187.020 284.620 187.660 ;
        RECT 0.270 185.660 284.620 187.020 ;
        RECT 0.270 183.580 287.435 185.660 ;
        RECT 4.400 181.580 284.620 183.580 ;
        RECT 0.270 179.500 287.435 181.580 ;
        RECT 4.400 178.140 287.435 179.500 ;
        RECT 4.400 177.500 284.620 178.140 ;
        RECT 0.270 176.140 284.620 177.500 ;
        RECT 0.270 175.420 287.435 176.140 ;
        RECT 4.400 174.060 287.435 175.420 ;
        RECT 4.400 173.420 284.620 174.060 ;
        RECT 0.270 172.060 284.620 173.420 ;
        RECT 0.270 169.980 287.435 172.060 ;
        RECT 4.400 168.620 287.435 169.980 ;
        RECT 4.400 167.980 284.620 168.620 ;
        RECT 0.270 166.620 284.620 167.980 ;
        RECT 0.270 165.900 287.435 166.620 ;
        RECT 4.400 164.540 287.435 165.900 ;
        RECT 4.400 163.900 284.620 164.540 ;
        RECT 0.270 162.540 284.620 163.900 ;
        RECT 0.270 160.460 287.435 162.540 ;
        RECT 4.400 158.460 284.620 160.460 ;
        RECT 0.270 156.380 287.435 158.460 ;
        RECT 4.400 155.020 287.435 156.380 ;
        RECT 4.400 154.380 284.620 155.020 ;
        RECT 0.270 153.020 284.620 154.380 ;
        RECT 0.270 152.300 287.435 153.020 ;
        RECT 4.400 150.940 287.435 152.300 ;
        RECT 4.400 150.300 284.620 150.940 ;
        RECT 0.270 148.940 284.620 150.300 ;
        RECT 0.270 146.860 287.435 148.940 ;
        RECT 4.400 144.860 284.620 146.860 ;
        RECT 0.270 142.780 287.435 144.860 ;
        RECT 4.400 141.420 287.435 142.780 ;
        RECT 4.400 140.780 284.620 141.420 ;
        RECT 0.270 139.420 284.620 140.780 ;
        RECT 0.270 138.700 287.435 139.420 ;
        RECT 4.400 137.340 287.435 138.700 ;
        RECT 4.400 136.700 284.620 137.340 ;
        RECT 0.270 135.340 284.620 136.700 ;
        RECT 0.270 133.260 287.435 135.340 ;
        RECT 4.400 131.260 284.620 133.260 ;
        RECT 0.270 129.180 287.435 131.260 ;
        RECT 4.400 127.820 287.435 129.180 ;
        RECT 4.400 127.180 284.620 127.820 ;
        RECT 0.270 125.820 284.620 127.180 ;
        RECT 0.270 123.740 287.435 125.820 ;
        RECT 4.400 121.740 284.620 123.740 ;
        RECT 0.270 119.660 287.435 121.740 ;
        RECT 4.400 118.300 287.435 119.660 ;
        RECT 4.400 117.660 284.620 118.300 ;
        RECT 0.270 116.300 284.620 117.660 ;
        RECT 0.270 115.580 287.435 116.300 ;
        RECT 4.400 114.220 287.435 115.580 ;
        RECT 4.400 113.580 284.620 114.220 ;
        RECT 0.270 112.220 284.620 113.580 ;
        RECT 0.270 110.140 287.435 112.220 ;
        RECT 4.400 108.140 284.620 110.140 ;
        RECT 0.270 106.060 287.435 108.140 ;
        RECT 4.400 104.700 287.435 106.060 ;
        RECT 4.400 104.060 284.620 104.700 ;
        RECT 0.270 102.700 284.620 104.060 ;
        RECT 0.270 101.980 287.435 102.700 ;
        RECT 4.400 100.620 287.435 101.980 ;
        RECT 4.400 99.980 284.620 100.620 ;
        RECT 0.270 98.620 284.620 99.980 ;
        RECT 0.270 96.540 287.435 98.620 ;
        RECT 4.400 94.540 284.620 96.540 ;
        RECT 0.270 92.460 287.435 94.540 ;
        RECT 4.400 91.100 287.435 92.460 ;
        RECT 4.400 90.460 284.620 91.100 ;
        RECT 0.270 89.100 284.620 90.460 ;
        RECT 0.270 88.380 287.435 89.100 ;
        RECT 4.400 87.020 287.435 88.380 ;
        RECT 4.400 86.380 284.620 87.020 ;
        RECT 0.270 85.020 284.620 86.380 ;
        RECT 0.270 82.940 287.435 85.020 ;
        RECT 4.400 81.580 287.435 82.940 ;
        RECT 4.400 80.940 284.620 81.580 ;
        RECT 0.270 79.580 284.620 80.940 ;
        RECT 0.270 78.860 287.435 79.580 ;
        RECT 4.400 77.500 287.435 78.860 ;
        RECT 4.400 76.860 284.620 77.500 ;
        RECT 0.270 75.500 284.620 76.860 ;
        RECT 0.270 73.420 287.435 75.500 ;
        RECT 4.400 71.420 284.620 73.420 ;
        RECT 0.270 69.340 287.435 71.420 ;
        RECT 4.400 67.980 287.435 69.340 ;
        RECT 4.400 67.340 284.620 67.980 ;
        RECT 0.270 65.980 284.620 67.340 ;
        RECT 0.270 65.260 287.435 65.980 ;
        RECT 4.400 63.900 287.435 65.260 ;
        RECT 4.400 63.260 284.620 63.900 ;
        RECT 0.270 61.900 284.620 63.260 ;
        RECT 0.270 59.820 287.435 61.900 ;
        RECT 4.400 57.820 284.620 59.820 ;
        RECT 0.270 55.740 287.435 57.820 ;
        RECT 4.400 54.380 287.435 55.740 ;
        RECT 4.400 53.740 284.620 54.380 ;
        RECT 0.270 52.380 284.620 53.740 ;
        RECT 0.270 51.660 287.435 52.380 ;
        RECT 4.400 50.300 287.435 51.660 ;
        RECT 4.400 49.660 284.620 50.300 ;
        RECT 0.270 48.300 284.620 49.660 ;
        RECT 0.270 46.220 287.435 48.300 ;
        RECT 4.400 44.220 284.620 46.220 ;
        RECT 0.270 42.140 287.435 44.220 ;
        RECT 4.400 40.780 287.435 42.140 ;
        RECT 4.400 40.140 284.620 40.780 ;
        RECT 0.270 38.780 284.620 40.140 ;
        RECT 0.270 36.700 287.435 38.780 ;
        RECT 4.400 34.700 284.620 36.700 ;
        RECT 0.270 32.620 287.435 34.700 ;
        RECT 4.400 31.260 287.435 32.620 ;
        RECT 4.400 30.620 284.620 31.260 ;
        RECT 0.270 29.260 284.620 30.620 ;
        RECT 0.270 28.540 287.435 29.260 ;
        RECT 4.400 27.180 287.435 28.540 ;
        RECT 4.400 26.540 284.620 27.180 ;
        RECT 0.270 25.180 284.620 26.540 ;
        RECT 0.270 23.100 287.435 25.180 ;
        RECT 4.400 21.100 284.620 23.100 ;
        RECT 0.270 19.020 287.435 21.100 ;
        RECT 4.400 17.660 287.435 19.020 ;
        RECT 4.400 17.020 284.620 17.660 ;
        RECT 0.270 15.660 284.620 17.020 ;
        RECT 0.270 14.940 287.435 15.660 ;
        RECT 4.400 13.580 287.435 14.940 ;
        RECT 4.400 12.940 284.620 13.580 ;
        RECT 0.270 11.580 284.620 12.940 ;
        RECT 0.270 9.500 287.435 11.580 ;
        RECT 4.400 7.500 284.620 9.500 ;
        RECT 0.270 5.420 287.435 7.500 ;
        RECT 4.400 4.060 287.435 5.420 ;
        RECT 4.400 3.420 284.620 4.060 ;
        RECT 0.270 2.060 284.620 3.420 ;
        RECT 0.270 0.175 287.435 2.060 ;
      LAYER met4 ;
        RECT 0.295 288.960 272.945 294.265 ;
        RECT 0.295 10.240 20.640 288.960 ;
        RECT 23.040 10.240 97.440 288.960 ;
        RECT 99.840 10.240 174.240 288.960 ;
        RECT 176.640 10.240 251.040 288.960 ;
        RECT 253.440 10.240 272.945 288.960 ;
        RECT 0.295 0.855 272.945 10.240 ;
  END
END both
END LIBRARY

